* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph1p3_clk_part                               *
* Netlisted  : Wed Nov  6 19:52:05 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_3 D_drain_1 S_source_0 3 B
** N=5 EP=4 FDC=1
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.2573 scb=0.0194507 scc=0.000476441 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_4 S_source_0 D_drain_1 3 4
** N=4 EP=4 FDC=1
M0 D_drain_1 3 S_source_0 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_5                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_5 D_drain_1 S_source_0 3 B
** N=5 EP=4 FDC=1
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.7106 scb=0.0166317 scc=0.000311047 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part CLK D Out gnd! vdd!
** N=6 EP=5 FDC=4
X2 Out D CLK vdd! pmos1v_CDNS_3 $T=1890 2460 0 0 $X=1470 $Y=2260
X3 gnd! 2 CLK gnd! nmos1v_CDNS_4 $T=710 860 0 0 $X=290 $Y=660
X4 D Out 2 gnd! nmos1v_CDNS_4 $T=1890 860 0 0 $X=1470 $Y=660
X5 2 vdd! CLK vdd! pmos1v_CDNS_5 $T=710 2460 0 0 $X=290 $Y=2260
.ends ph1p3_clk_part
