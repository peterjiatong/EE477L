* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph3_sytolic_array                            *
* Netlisted  : Sun Dec  8 18:33:48 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_new                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_new vdd gnd 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 4 3 gnd gnd g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.3086 scb=0.00950139 scc=0.000267597 $X=1140 $Y=930 $dt=0
.ends INV_1X_new

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X_small                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X_small 1 vdd! gnd! 4 out
*.DEVICECLIMB
** N=6 EP=5 FDC=2
M0 6 1 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=810 $Y=1000 $dt=0
M1 out 4 6 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=2050 $Y=1000 $dt=0
.ends NAND2_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND in_A vdd! gnd! in_B out 6
*.DEVICECLIMB
** N=7 EP=6 FDC=3
X0 vdd! gnd! 6 out INV_1X_new $T=2480 -10 0 0 $X=2410 $Y=0
X1 in_A vdd! gnd! in_B 6 NAND2_1X_small $T=-110 -70 0 0 $X=10 $Y=0
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR_small                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR_small in_A vdd! gnd! in_B out 6 8
*.DEVICECLIMB
** N=10 EP=7 FDC=9
M0 8 in_A gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.45462 scb=0.00478425 scc=6.8709e-05 $X=700 $Y=590 $dt=0
M1 7 in_B gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=2110 $Y=580 $dt=0
M2 9 7 gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=3270 $Y=580 $dt=0
M3 out 8 9 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=4610 $Y=580 $dt=0
M4 10 in_B gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 $X=6140 $Y=600 $dt=0
M5 out in_A 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=7250 $Y=650 $dt=0
M6 7 in_B vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.1869 scb=0.0086398 scc=0.00051649 $X=2110 $Y=2170 $dt=1
M7 6 7 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3270 $Y=2160 $dt=1
M8 6 8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4610 $Y=2160 $dt=1
.ends XOR_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder inA gnd! vdd! inB S C 8 9 13
*.DEVICECLIMB
** N=13 EP=9 FDC=12
X6 inA vdd! gnd! inB C 9 AND $T=7790 0 0 0 $X=7800 $Y=0
X7 inA vdd! gnd! inB S 13 8 XOR_small $T=0 0 0 0 $X=0 $Y=0
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_1X_small                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_1X_small vdd! gnd! 3 4 5
*.DEVICECLIMB
** N=6 EP=5 FDC=2
M0 6 3 gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1000 $Y=830 $dt=0
M1 4 5 6 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1210 $Y=830 $dt=0
.ends NAND_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_2X_small1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_2X_small1 vdd! gnd! out 4 5
*.DEVICECLIMB
** N=6 EP=5 FDC=2
M0 6 4 gnd! gnd! g45n1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=7.66878 scb=0.00580736 scc=7.77234e-05 $X=940 $Y=890 $dt=0
M1 out 5 6 gnd! g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=11.676 scb=0.0124835 scc=0.000479408 $X=940 $Y=1100 $dt=0
.ends NAND_2X_small1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR1 vdd! gnd! 3 4 5 6 7 9
*.DEVICECLIMB
** N=10 EP=8 FDC=6
M0 6 3 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=830 $Y=840 $dt=0
M1 7 4 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1790 $Y=840 $dt=0
M2 8 4 gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=3120 $Y=780 $dt=0
M3 5 6 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4126 scb=0.0095497 scc=0.000351079 $X=4090 $Y=760 $dt=0
M4 gnd! 7 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=5050 $Y=770 $dt=0
M5 5 3 8 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=6010 $Y=770 $dt=0
.ends XOR1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder1_small                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder1_small inA vdd! inB gnd! Cin_ S Cout 8 9 10
+ 11 12 13 14 22 23
*.DEVICECLIMB
** N=23 EP=16 FDC=18
X26 vdd! gnd! inA 10 inB NAND_1X_small $T=16970 30 0 0 $X=16540 $Y=10
X27 vdd! gnd! 9 Cout 10 NAND_1X_small $T=19810 30 0 0 $X=19380 $Y=10
X28 vdd! gnd! 9 Cin_ 8 NAND_2X_small1 $T=13690 -10 0 0 $X=13700 $Y=10
X29 vdd! gnd! inA inB 8 11 12 22 XOR1 $T=-40 30 0 0 $X=20 $Y=10
X30 vdd! gnd! Cin_ 8 S 13 14 23 XOR1 $T=6800 30 0 0 $X=6860 $Y=10
.ends full_adder1_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: multiplier                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt multiplier a3 gnd! b0 b2 b3 vdd! a2 a1 b1 z6
+ a0 z7 z3 z0 z5 z4 z2 z1
** N=238 EP=18 FDC=456
X273 a3 vdd! gnd! b3 43 77 AND $T=40 14460 1 0 $X=50 $Y=10660
X274 a3 vdd! gnd! b2 21 76 AND $T=40 14420 0 0 $X=50 $Y=14420
X275 a3 vdd! gnd! b0 20 75 AND $T=40 21740 0 0 $X=50 $Y=21740
X276 a2 vdd! gnd! b3 39 80 AND $T=4440 14460 1 0 $X=4450 $Y=10660
X277 a2 vdd! gnd! b2 24 79 AND $T=4440 14420 0 0 $X=4450 $Y=14420
X278 a3 vdd! gnd! b1 23 78 AND $T=4440 21740 0 0 $X=4450 $Y=21740
X279 a1 vdd! gnd! b3 38 83 AND $T=8840 14460 1 0 $X=8850 $Y=10660
X280 a1 vdd! gnd! b2 26 82 AND $T=8840 14420 0 0 $X=8850 $Y=14420
X281 b0 vdd! gnd! a2 35 81 AND $T=8840 21740 0 0 $X=8850 $Y=21740
X282 a0 vdd! gnd! b3 50 93 AND $T=13240 14460 1 0 $X=13250 $Y=10660
X283 a0 vdd! gnd! b2 45 92 AND $T=13240 14420 0 0 $X=13250 $Y=14420
X284 b1 vdd! gnd! a2 27 91 AND $T=13240 21740 0 0 $X=13250 $Y=21740
X285 b0 vdd! gnd! a1 30 104 AND $T=17880 21740 0 0 $X=17890 $Y=21740
X286 b1 vdd! gnd! a1 33 126 AND $T=22280 21740 0 0 $X=22290 $Y=21740
X287 b0 vdd! gnd! a0 z0 127 AND $T=26680 21740 0 0 $X=26690 $Y=21740
X288 b1 vdd! gnd! a0 31 131 AND $T=31080 21740 0 0 $X=31090 $Y=21740
X289 23 gnd! vdd! 37 22 25 73 74 225 half_adder $T=50 21780 1 0 $X=50 $Y=17980
X290 50 gnd! vdd! 48 z3 46 102 103 228 half_adder $T=17640 14460 1 0 $X=17640 $Y=10660
X291 45 gnd! vdd! 47 z2 49 129 130 237 half_adder $T=29830 14460 1 0 $X=29830 $Y=10660
X292 30 gnd! vdd! 31 z1 32 133 134 238 half_adder $T=34210 21780 1 0 $X=34210 $Y=17980
X293 22 vdd! 24 gnd! 28 36 19 67 70 71
+ 65 66 68 69 223 224 full_adder1_small $T=22270 7090 1 180 $X=20 $Y=7100
X294 43 vdd! 34 gnd! 29 z6 z7 60 63 64
+ 58 59 61 62 221 222 full_adder1_small $T=30 -230 0 0 $X=50 $Y=-220
X295 21 vdd! 25 gnd! 19 44 34 53 56 57
+ 51 52 54 55 219 220 full_adder1_small $T=30 7150 1 0 $X=50 $Y=3340
X296 20 vdd! 27 gnd! 41 40 37 86 89 90
+ 84 85 87 88 226 227 full_adder1_small $T=12230 21790 1 0 $X=12250 $Y=17980
X297 33 vdd! 35 gnd! 32 47 41 96 99 100
+ 94 95 97 98 229 230 full_adder1_small $T=17850 14410 0 0 $X=17870 $Y=14420
X298 39 vdd! 44 gnd! 42 z5 29 121 124 125
+ 119 120 122 123 235 236 full_adder1_small $T=21990 -230 0 0 $X=22010 $Y=-220
X299 38 vdd! 36 gnd! 46 z4 42 114 117 118
+ 112 113 115 116 233 234 full_adder1_small $T=21990 7150 1 0 $X=22010 $Y=3340
X300 26 vdd! 40 gnd! 49 48 28 107 110 111
+ 105 106 108 109 231 232 full_adder1_small $T=21990 7090 0 0 $X=22010 $Y=7100
M0 77 a3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=11610 $dt=1
M1 76 a3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=16790 $dt=1
M2 75 a3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=24110 $dt=1
M3 73 23 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=16.2188 scb=0.0173423 scc=0.000698846 $X=750 $Y=18640 $dt=1
M4 58 43 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=2120 $dt=1
M5 51 21 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=4320 $dt=1
M6 19 71 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=1070 $Y=9450 $dt=1
M7 vdd! 70 19 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=1480 $Y=9450 $dt=1
M8 59 34 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=2120 $dt=1
M9 52 25 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=4320 $dt=1
M10 77 b3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=11600 $dt=1
M11 76 b2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=16800 $dt=1
M12 75 b0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=24120 $dt=1
M13 221 34 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=1880 $dt=1
M14 219 25 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=4080 $dt=1
M15 43 77 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=11580 $dt=1
M16 21 76 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=16820 $dt=1
M17 20 75 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=24140 $dt=1
M18 71 24 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=3910 $Y=9450 $dt=1
M19 60 58 221 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=1940 $dt=1
M20 53 51 219 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=4020 $dt=1
M21 vdd! 22 71 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=4320 $Y=9450 $dt=1
M22 60 59 221 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=1940 $dt=1
M23 53 52 219 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=4020 $dt=1
M24 80 a2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=11610 $dt=1
M25 79 a2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=16790 $dt=1
M26 78 a3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=24110 $dt=1
M27 221 43 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=1940 $dt=1
M28 219 21 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=4020 $dt=1
M29 22 37 225 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=6190 $Y=18700 $dt=1
M30 80 b3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=11600 $dt=1
M31 79 b2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=16800 $dt=1
M32 78 b1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=24120 $dt=1
M33 70 67 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=6890 $Y=9230 $dt=1
M34 vdd! 28 70 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=7300 $Y=9230 $dt=1
M35 22 23 225 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=7300 $Y=18660 $dt=1
M36 61 29 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=2120 $dt=1
M37 54 19 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=4320 $dt=1
M38 39 80 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=11580 $dt=1
M39 24 79 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=16820 $dt=1
M40 23 78 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=24140 $dt=1
M41 74 23 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=8540 $Y=18930 $dt=1
M42 62 60 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=2120 $dt=1
M43 55 53 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=4320 $dt=1
M44 vdd! 28 224 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=9370 $Y=9260 $dt=1
M45 83 a1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=11610 $dt=1
M46 82 a1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=16790 $dt=1
M47 81 b0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=24110 $dt=1
M48 74 37 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=9780 $Y=18920 $dt=1
M49 222 60 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=1880 $dt=1
M50 220 53 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=4080 $dt=1
M51 224 69 36 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10330 $Y=9260 $dt=1
M52 83 b3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=11600 $dt=1
M53 82 b2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=16800 $dt=1
M54 81 a2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=24120 $dt=1
M55 z6 61 222 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=1940 $dt=1
M56 44 54 220 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=4020 $dt=1
M57 224 68 36 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11290 $Y=9260 $dt=1
M58 25 74 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=11460 $Y=18900 $dt=1
M59 z6 62 222 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=1940 $dt=1
M60 44 55 220 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=4020 $dt=1
M61 vdd! 67 224 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=12260 $Y=9200 $dt=1
M62 38 83 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=11580 $dt=1
M63 26 82 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=16820 $dt=1
M64 35 81 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=24140 $dt=1
M65 222 29 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=1940 $dt=1
M66 220 19 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=4020 $dt=1
M67 84 20 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13020 $Y=18960 $dt=1
M68 vdd! 67 69 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13590 $Y=9440 $dt=1
M69 93 a0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=11610 $dt=1
M70 92 a0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=16790 $dt=1
M71 91 b1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=24110 $dt=1
M72 85 27 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13980 $Y=18960 $dt=1
M73 vdd! 28 68 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=14550 $Y=9440 $dt=1
M74 63 29 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=1910 $dt=1
M75 56 19 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=4050 $dt=1
M76 93 b3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=11600 $dt=1
M77 92 b2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=16800 $dt=1
M78 91 a2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=24120 $dt=1
M79 226 27 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=15310 $Y=18720 $dt=1
M80 vdd! 60 63 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=1910 $dt=1
M81 vdd! 53 56 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=4050 $dt=1
M82 vdd! 22 223 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16210 $Y=9260 $dt=1
M83 86 84 226 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16280 $Y=18660 $dt=1
M84 50 93 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=11580 $dt=1
M85 45 92 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=16820 $dt=1
M86 27 91 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=24140 $dt=1
M87 223 66 67 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17170 $Y=9260 $dt=1
M88 86 85 226 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17240 $Y=18660 $dt=1
M89 64 43 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=2130 $dt=1
M90 57 21 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=4310 $dt=1
M91 223 65 67 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18130 $Y=9260 $dt=1
M92 226 20 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18200 $Y=18660 $dt=1
M93 vdd! 34 64 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=2130 $dt=1
M94 vdd! 25 57 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=4310 $dt=1
M95 102 50 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=18340 $Y=11320 $dt=1
M96 104 b0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=18580 $Y=24110 $dt=1
M97 94 33 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=18640 $Y=16760 $dt=1
M98 vdd! 24 223 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=19100 $Y=9200 $dt=1
M99 95 35 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19600 $Y=16760 $dt=1
M100 104 a1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=19820 $Y=24120 $dt=1
M101 87 41 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19860 $Y=18960 $dt=1
M102 vdd! 24 66 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20430 $Y=9440 $dt=1
M103 z7 63 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=2130 $dt=1
M104 34 56 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=4310 $dt=1
M105 88 86 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20820 $Y=18960 $dt=1
M106 229 35 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=20930 $Y=16520 $dt=1
M107 vdd! 64 z7 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=2130 $dt=1
M108 vdd! 57 34 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=4310 $dt=1
M109 vdd! 22 65 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=21390 $Y=9440 $dt=1
M110 30 104 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=21500 $Y=24140 $dt=1
M111 96 94 229 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=21900 $Y=16580 $dt=1
M112 227 86 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=22150 $Y=18720 $dt=1
M113 119 39 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=2120 $dt=1
M114 112 38 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=4320 $dt=1
M115 105 26 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=9440 $dt=1
M116 96 95 229 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=22860 $Y=16580 $dt=1
M117 126 b1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=22980 $Y=24110 $dt=1
M118 40 87 227 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23120 $Y=18660 $dt=1
M119 120 44 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=2120 $dt=1
M120 113 36 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=4320 $dt=1
M121 106 40 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=9440 $dt=1
M122 z3 48 228 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=23780 $Y=11380 $dt=1
M123 229 33 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23820 $Y=16580 $dt=1
M124 40 88 227 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24080 $Y=18660 $dt=1
M125 126 a1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=24220 $Y=24120 $dt=1
M126 z3 50 228 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24890 $Y=11340 $dt=1
M127 227 41 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=25040 $Y=18660 $dt=1
M128 235 44 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=1880 $dt=1
M129 233 36 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=4080 $dt=1
M130 231 40 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=9200 $dt=1
M131 97 32 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=25480 $Y=16760 $dt=1
M132 33 126 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=25900 $Y=24140 $dt=1
M133 121 119 235 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=1940 $dt=1
M134 114 112 233 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=4020 $dt=1
M135 107 105 231 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=9260 $dt=1
M136 103 50 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26130 $Y=11610 $dt=1
M137 98 96 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=26440 $Y=16760 $dt=1
M138 121 120 235 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=1940 $dt=1
M139 114 113 233 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=4020 $dt=1
M140 107 106 231 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=9260 $dt=1
M141 89 41 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27110 $Y=18690 $dt=1
M142 103 48 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27370 $Y=11600 $dt=1
M143 127 b0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=27380 $Y=24110 $dt=1
M144 vdd! 86 89 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27520 $Y=18690 $dt=1
M145 230 96 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=27770 $Y=16520 $dt=1
M146 235 39 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=1940 $dt=1
M147 233 38 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=4020 $dt=1
M148 231 26 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=9260 $dt=1
M149 127 a0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=28620 $Y=24120 $dt=1
M150 47 97 230 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28740 $Y=16580 $dt=1
M151 46 103 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=29050 $Y=11580 $dt=1
M152 122 42 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=2120 $dt=1
M153 115 46 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=4320 $dt=1
M154 108 49 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=9440 $dt=1
M155 47 98 230 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=29700 $Y=16580 $dt=1
M156 90 20 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30090 $Y=18950 $dt=1
M157 z0 127 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=30300 $Y=24140 $dt=1
M158 vdd! 27 90 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30500 $Y=18950 $dt=1
M159 129 45 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=30530 $Y=11320 $dt=1
M160 123 121 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=2120 $dt=1
M161 116 114 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=4320 $dt=1
M162 109 107 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=9440 $dt=1
M163 230 32 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=30660 $Y=16580 $dt=1
M164 131 b1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=31780 $Y=24110 $dt=1
M165 236 121 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=1880 $dt=1
M166 234 114 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=4080 $dt=1
M167 232 107 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=9200 $dt=1
M168 99 32 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=32730 $Y=16550 $dt=1
M169 z5 122 236 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=1940 $dt=1
M170 z4 115 234 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=4020 $dt=1
M171 48 108 232 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=9260 $dt=1
M172 37 89 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=32930 $Y=18950 $dt=1
M173 131 a0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=33020 $Y=24120 $dt=1
M174 vdd! 96 99 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=33140 $Y=16550 $dt=1
M175 vdd! 90 37 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=33340 $Y=18950 $dt=1
M176 z5 123 236 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=1940 $dt=1
M177 z4 116 234 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=4020 $dt=1
M178 48 109 232 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=9260 $dt=1
M179 31 131 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=34700 $Y=24140 $dt=1
M180 236 42 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=1940 $dt=1
M181 234 46 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=4020 $dt=1
M182 232 49 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=9260 $dt=1
M183 133 30 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=34910 $Y=18640 $dt=1
M184 100 33 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=35710 $Y=16770 $dt=1
M185 z2 47 237 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=35970 $Y=11380 $dt=1
M186 vdd! 35 100 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=36120 $Y=16770 $dt=1
M187 124 42 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=1910 $dt=1
M188 117 46 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=4050 $dt=1
M189 110 49 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=9230 $dt=1
M190 z2 45 237 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=37080 $Y=11340 $dt=1
M191 vdd! 121 124 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=1910 $dt=1
M192 vdd! 114 117 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=4050 $dt=1
M193 vdd! 107 110 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=9230 $dt=1
M194 130 45 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=38320 $Y=11610 $dt=1
M195 41 99 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=38550 $Y=16770 $dt=1
M196 vdd! 100 41 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=38960 $Y=16770 $dt=1
M197 130 47 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=39560 $Y=11600 $dt=1
M198 125 39 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=2130 $dt=1
M199 118 38 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=4310 $dt=1
M200 111 26 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=9450 $dt=1
M201 vdd! 44 125 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=2130 $dt=1
M202 vdd! 36 118 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=4310 $dt=1
M203 vdd! 40 111 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=9450 $dt=1
M204 z1 31 238 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.2705 scb=0.0126902 scc=0.000796523 $X=40350 $Y=18700 $dt=1
M205 49 130 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=41240 $Y=11580 $dt=1
M206 z1 30 238 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=41460 $Y=18660 $dt=1
M207 29 124 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=2130 $dt=1
M208 42 117 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=4310 $dt=1
M209 28 110 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=42690 $Y=9450 $dt=1
M210 134 30 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42700 $Y=18930 $dt=1
M211 vdd! 125 29 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=2130 $dt=1
M212 vdd! 118 42 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=4310 $dt=1
M213 vdd! 111 28 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=43100 $Y=9450 $dt=1
M214 134 31 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43940 $Y=18920 $dt=1
M215 32 134 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=45620 $Y=18900 $dt=1
.ends multiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_43                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_43 2 3 5 6 8
*.DEVICECLIMB
** N=14 EP=5 FDC=2
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=810 $Y=710 $dt=0
M1 8 6 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=4640 $Y=580 $dt=0
.ends cellTmpl_CDNS_43

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X S A vdd! gnd! B out
** N=12 EP=6 FDC=12
X20 gnd! S 7 8 out cellTmpl_CDNS_43 $T=-60 -5080 0 0 $X=-180 $Y=-5220
M0 9 A 8 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1780 $Y=-4420 $dt=0
M1 gnd! 7 9 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1990 $Y=-4420 $dt=0
M2 10 S gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3160 $Y=-4430 $dt=0
M3 8 B 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3370 $Y=-4430 $dt=0
M4 7 S vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=750 $Y=-2850 $dt=1
M5 11 A 8 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1780 $Y=-3120 $dt=1
M6 vdd! S 11 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1990 $Y=-3120 $dt=1
M7 12 7 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3160 $Y=-3190 $dt=1
M8 8 B 12 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3370 $Y=-3190 $dt=1
M9 out 8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.2373 scb=0.0194294 scc=0.00149528 $X=4580 $Y=-3180 $dt=1
.ends MUX_2to1___2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FA_4bit                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FA_4bit B0 B1 B2 B3 vdd! A0 gnd! A1 A2 A3
+ Cin_rrr S0 S1 S2 S3 Cout3
** N=83 EP=16 FDC=144
X21 A0 vdd! B0 gnd! Cin_rrr S0 18 43 46 47
+ 41 42 44 45 82 83 full_adder1_small $T=-90 -130 0 0 $X=-70 $Y=-120
X22 A1 vdd! B1 gnd! 18 S1 17 36 39 40
+ 34 35 37 38 80 81 full_adder1_small $T=-90 7250 1 0 $X=-70 $Y=3440
X23 A2 vdd! B2 gnd! 17 S2 19 29 32 33
+ 27 28 30 31 78 79 full_adder1_small $T=-90 7190 0 0 $X=-70 $Y=7200
X24 A3 vdd! B3 gnd! 19 S3 Cout3 22 25 26
+ 20 21 23 24 76 77 full_adder1_small $T=-90 14570 1 0 $X=-70 $Y=10760
M0 41 A0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=2220 $dt=1
M1 34 A1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=4420 $dt=1
M2 27 A2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=9540 $dt=1
M3 20 A3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=11740 $dt=1
M4 42 B0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=2220 $dt=1
M5 35 B1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=4420 $dt=1
M6 28 B2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=9540 $dt=1
M7 21 B3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=11740 $dt=1
M8 82 B0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=1980 $dt=1
M9 80 B1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=4180 $dt=1
M10 78 B2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=9300 $dt=1
M11 76 B3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=11500 $dt=1
M12 43 41 82 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=2040 $dt=1
M13 36 34 80 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=4120 $dt=1
M14 29 27 78 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=9360 $dt=1
M15 22 20 76 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=11440 $dt=1
M16 43 42 82 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=2040 $dt=1
M17 36 35 80 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=4120 $dt=1
M18 29 28 78 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=9360 $dt=1
M19 22 21 76 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=11440 $dt=1
M20 82 A0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=2040 $dt=1
M21 80 A1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=4120 $dt=1
M22 78 A2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=9360 $dt=1
M23 76 A3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=11440 $dt=1
M24 44 Cin_rrr vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=2220 $dt=1
M25 37 18 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=4420 $dt=1
M26 30 17 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=9540 $dt=1
M27 23 19 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=11740 $dt=1
M28 45 43 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=2220 $dt=1
M29 38 36 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=4420 $dt=1
M30 31 29 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=9540 $dt=1
M31 24 22 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=11740 $dt=1
M32 83 43 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=1980 $dt=1
M33 81 36 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=4180 $dt=1
M34 79 29 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=9300 $dt=1
M35 77 22 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=11500 $dt=1
M36 S0 44 83 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=2040 $dt=1
M37 S1 37 81 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=4120 $dt=1
M38 S2 30 79 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=9360 $dt=1
M39 S3 23 77 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=11440 $dt=1
M40 S0 45 83 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=2040 $dt=1
M41 S1 38 81 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=4120 $dt=1
M42 S2 31 79 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=9360 $dt=1
M43 S3 24 77 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=11440 $dt=1
M44 83 Cin_rrr vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=2040 $dt=1
M45 81 18 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=4120 $dt=1
M46 79 17 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=9360 $dt=1
M47 77 19 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=11440 $dt=1
M48 46 Cin_rrr vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=2010 $dt=1
M49 39 18 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=4150 $dt=1
M50 32 17 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=9330 $dt=1
M51 25 19 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=11470 $dt=1
M52 vdd! 43 46 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=2010 $dt=1
M53 vdd! 36 39 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=4150 $dt=1
M54 vdd! 29 32 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=9330 $dt=1
M55 vdd! 22 25 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=11470 $dt=1
M56 47 A0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=2230 $dt=1
M57 40 A1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=4410 $dt=1
M58 33 A2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=9550 $dt=1
M59 26 A3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=11730 $dt=1
M60 vdd! B0 47 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=2230 $dt=1
M61 vdd! B1 40 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=4410 $dt=1
M62 vdd! B2 33 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=9550 $dt=1
M63 vdd! B3 26 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=11730 $dt=1
M64 18 46 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=2230 $dt=1
M65 17 39 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=4410 $dt=1
M66 19 32 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=9550 $dt=1
M67 Cout3 25 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=11730 $dt=1
M68 vdd! 47 18 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=2230 $dt=1
M69 vdd! 40 17 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=4410 $dt=1
M70 vdd! 33 19 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=9550 $dt=1
M71 vdd! 26 Cout3 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=11730 $dt=1
.ends FA_4bit

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small in vdd! gnd! out
** N=4 EP=4 FDC=2
M0 out in gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7353 scb=0.0117274 scc=0.000445561 $X=1070 $Y=980 $dt=0
M1 out in vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8675 scb=0.0146094 scc=0.000688105 $X=1070 $Y=2220 $dt=1
.ends INV_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 10badder                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 10badder in_A_8 Cin vdd! gnd! in_B_8 in_A_4 in_A_0 in_B_7 in_B_6 in_B_5
+ in_B_3 in_B_2 in_B_1 in_B_0 in_A_1 in_A_2 in_A_3 in_B_4 in_A_5 in_A_6
+ in_A_7 S8 in_B_9 in_A_9 S0 S3 S2 S1 S7 S6
+ S5 S4 S9 Cout 50 51 64 65 66 67
+ 68 69 70 149 150 151 152 153 154 155
+ 256 257 266 267
*.DEVICECLIMB
** N=267 EP=54 FDC=483
X148 vdd! gnd! 40 56 42 NAND_1X_small $T=53960 20720 0 0 $X=53530 $Y=20700
X149 vdd! gnd! 36 58 52 NAND_1X_small $T=55940 28040 0 180 $X=53530 $Y=24260
X150 vdd! gnd! 38 54 44 NAND_1X_small $T=53960 28040 0 0 $X=53530 $Y=28020
X151 vdd! gnd! 41 57 43 NAND_1X_small $T=53960 35360 0 0 $X=53530 $Y=35340
X152 vdd! gnd! 37 59 53 NAND_1X_small $T=55940 42680 0 180 $X=53530 $Y=38900
X153 vdd! gnd! 39 55 45 NAND_1X_small $T=53960 42680 0 0 $X=53530 $Y=42660
X154 vdd! gnd! in_B_0 in_A_0 42 85 86 265 XOR1 $T=56070 20720 0 0 $X=56130 $Y=20700
X155 vdd! gnd! in_A_1 in_B_1 40 83 84 264 XOR1 $T=56070 28040 1 0 $X=56130 $Y=24260
X156 vdd! gnd! in_A_2 in_B_2 44 81 82 263 XOR1 $T=56070 28040 0 0 $X=56130 $Y=28020
X157 vdd! gnd! in_A_3 in_B_3 38 79 80 262 XOR1 $T=56070 35360 1 0 $X=56130 $Y=31580
X158 vdd! gnd! in_B_4 in_A_4 43 77 78 261 XOR1 $T=56070 35360 0 0 $X=56130 $Y=35340
X159 vdd! gnd! in_A_5 in_B_5 41 75 76 260 XOR1 $T=56070 42680 1 0 $X=56130 $Y=38900
X160 vdd! gnd! in_A_6 in_B_6 45 73 74 259 XOR1 $T=56070 42680 0 0 $X=56130 $Y=42660
X161 vdd! gnd! in_A_7 in_B_7 39 71 72 258 XOR1 $T=56070 50000 1 0 $X=56130 $Y=46220
X162 in_B_8 vdd! in_A_8 gnd! 50 S8 51 66 69 70
+ 64 65 67 68 256 257 full_adder1_small $T=50650 49970 0 0 $X=50670 $Y=49980
X163 in_A_9 vdd! in_B_9 gnd! 51 S9 Cout 151 154 155
+ 149 150 152 153 266 267 full_adder1_small $T=72610 49970 0 0 $X=72630 $Y=49980
X164 46 48 vdd! gnd! Cin 35 MUX_2to1___2X $T=56190 30160 0 180 $X=50640 $Y=31580
X165 47 49 vdd! gnd! 35 50 MUX_2to1___2X $T=56190 44800 0 180 $X=50640 $Y=46220
X166 in_B_0 in_B_1 in_B_2 in_B_3 vdd! in_A_0 gnd! in_A_1 in_A_2 in_A_3
+ Cin S0 S1 S2 S3 48 FA_4bit $T=64900 20820 0 0 $X=64250 $Y=20700
X167 in_B_4 in_B_5 in_B_6 in_B_7 vdd! in_A_4 gnd! in_A_5 in_A_6 in_A_7
+ 35 S4 S5 S6 S7 49 FA_4bit $T=64900 35460 0 0 $X=64250 $Y=35340
X168 56 vdd! gnd! 52 INV_1X_small $T=51530 20700 0 0 $X=51530 $Y=20700
X169 58 vdd! gnd! 46 INV_1X_small $T=51530 28060 1 0 $X=51530 $Y=24260
X170 54 vdd! gnd! 36 INV_1X_small $T=51530 28020 0 0 $X=51530 $Y=28020
X171 57 vdd! gnd! 53 INV_1X_small $T=51530 35340 0 0 $X=51530 $Y=35340
X172 59 vdd! gnd! 47 INV_1X_small $T=51530 42700 1 0 $X=51530 $Y=38900
X173 55 vdd! gnd! 37 INV_1X_small $T=51530 42660 0 0 $X=51530 $Y=42660
M0 64 in_B_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6612 scb=0.0167915 scc=0.000377457 $X=51440 $Y=52320 $dt=1
M1 58 52 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=25230 $dt=1
M2 59 53 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=39870 $dt=1
M3 56 40 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=23050 $dt=1
M4 54 38 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=30370 $dt=1
M5 57 41 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=37690 $dt=1
M6 55 39 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=45010 $dt=1
M7 vdd! 36 58 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=25230 $dt=1
M8 vdd! 37 59 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=39870 $dt=1
M9 vdd! 42 56 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=23050 $dt=1
M10 vdd! 44 54 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=30370 $dt=1
M11 vdd! 43 57 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=37690 $dt=1
M12 vdd! 45 55 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=45010 $dt=1
M13 85 in_B_0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=23040 $dt=1
M14 83 in_A_1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=25240 $dt=1
M15 81 in_A_2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=30360 $dt=1
M16 79 in_A_3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=32560 $dt=1
M17 77 in_B_4 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=37680 $dt=1
M18 75 in_A_5 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=39880 $dt=1
M19 73 in_A_6 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=45000 $dt=1
M20 71 in_A_7 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=47200 $dt=1
M21 86 in_A_0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=23040 $dt=1
M22 84 in_B_1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=25240 $dt=1
M23 82 in_B_2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=30360 $dt=1
M24 80 in_B_3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=32560 $dt=1
M25 78 in_A_4 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=37680 $dt=1
M26 76 in_B_5 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=39880 $dt=1
M27 74 in_B_6 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=45000 $dt=1
M28 72 in_B_7 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=47200 $dt=1
M29 265 in_A_0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=22800 $dt=1
M30 264 in_B_1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=25000 $dt=1
M31 263 in_B_2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=30120 $dt=1
M32 262 in_B_3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=32320 $dt=1
M33 261 in_A_4 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=37440 $dt=1
M34 260 in_B_5 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=39640 $dt=1
M35 259 in_B_6 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=44760 $dt=1
M36 258 in_B_7 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=46960 $dt=1
M37 42 85 265 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=22860 $dt=1
M38 40 83 264 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=24940 $dt=1
M39 44 81 263 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=30180 $dt=1
M40 38 79 262 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=32260 $dt=1
M41 43 77 261 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=37500 $dt=1
M42 41 75 260 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=39580 $dt=1
M43 45 73 259 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=44820 $dt=1
M44 39 71 258 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=46900 $dt=1
M45 42 86 265 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=22860 $dt=1
M46 40 84 264 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=24940 $dt=1
M47 44 82 263 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=30180 $dt=1
M48 38 80 262 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=32260 $dt=1
M49 43 78 261 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=37500 $dt=1
M50 41 76 260 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=39580 $dt=1
M51 45 74 259 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=44820 $dt=1
M52 39 72 258 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=46900 $dt=1
M53 265 in_B_0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=22860 $dt=1
M54 264 in_A_1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=24940 $dt=1
M55 263 in_A_2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=30180 $dt=1
M56 262 in_A_3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=32260 $dt=1
M57 261 in_B_4 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=37500 $dt=1
M58 260 in_A_5 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=39580 $dt=1
M59 259 in_A_6 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=44820 $dt=1
M60 258 in_A_7 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=46900 $dt=1
M61 Cout 154 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=93310 $Y=52330 $dt=1
M62 vdd! 155 Cout vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=93720 $Y=52330 $dt=1
.ends 10badder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_46                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_46 2 3 5
*.DEVICECLIMB
** N=5 EP=3 FDC=1
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=660 $Y=760 $dt=0
.ends cellTmpl_CDNS_46

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout in vdd! gnd! out
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X1 gnd! in out cellTmpl_CDNS_46 $T=120 140 0 0 $X=0 $Y=0
.ends INV_1X_small_layout

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part CLK vdd! gnd! D Out 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
M0 6 CLK gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=710 $Y=860 $dt=0
M1 Out 6 D gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1890 $Y=860 $dt=0
.ends ph1p3_clk_part

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_MSDFF                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_MSDFF vdd! CLK gnd! RST D Q 7 8 9 10
+ 11 12 13 14 15 16 17
*.DEVICECLIMB
** N=18 EP=17 FDC=15
X33 8 vdd! gnd! 10 12 NAND2_1X_small $T=3680 -70 0 0 $X=3800 $Y=0
X34 RST vdd! gnd! 10 INV_1X_small_layout $T=0 40 1 0 $X=0 $Y=-3760
X35 CLK vdd! gnd! 7 INV_1X_small_layout $T=0 0 0 0 $X=0 $Y=0
X36 Q vdd! gnd! 11 INV_1X_small_layout $T=4800 40 1 0 $X=4800 $Y=-3760
X37 12 vdd! gnd! 13 INV_1X_small_layout $T=6200 0 0 0 $X=6200 $Y=0
X38 9 vdd! gnd! Q INV_1X_small_layout $T=8600 40 1 0 $X=8600 $Y=-3760
X39 CLK vdd! gnd! D 8 14 ph1p3_clk_part $T=1400 0 0 0 $X=1400 $Y=0
X40 CLK vdd! gnd! 11 9 15 ph1p3_clk_part $T=2400 40 1 0 $X=2400 $Y=-3760
X41 7 vdd! gnd! 12 9 16 ph1p3_clk_part $T=6200 40 1 0 $X=6200 $Y=-3760
X42 7 vdd! gnd! 13 8 17 ph1p3_clk_part $T=7600 0 0 0 $X=7600 $Y=0
.ends ph1p3_MSDFF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X_ph2p2                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X_ph2p2 S A vdd! gnd! B out 7 8 11 12
*.DEVICECLIMB
** N=12 EP=10 FDC=6
X20 gnd! S 7 8 out cellTmpl_CDNS_43 $T=120 140 0 0 $X=0 $Y=0
M0 9 A 8 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1960 $Y=800 $dt=0
M1 gnd! 7 9 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=2170 $Y=800 $dt=0
M2 10 S gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3340 $Y=790 $dt=0
M3 8 B 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3550 $Y=790 $dt=0
.ends MUX_2to1___2X_ph2p2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p2_processing_element                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p2_processing_element A3 B0 B2 B3 gnd! RST CLK Cin A8 vdd!
+ B1 A_reg3 B_reg0 A1 A2 A0 B_reg1 A_reg2 A9 B_reg2
+ A_reg1 A_reg0 B_reg3 Sel Sel_reg Sum_out5 Sum_out0 Sum_out3 Sum_out9 Sum_out1
+ Sum_out8 Sum_out4 Sum_out2 Sum_out6 Sum_out7 Sum_in6 Sum_in9 Sum_in5 Sum_in8 Sum_in4
+ Sum_in7 Sum_in3 Sum_in2 Sum_in1 Sum_in0 63 64 69 70 75
+ 77 78 79 81 83 108 113 130 139 140
+ 141 158 159 176 185 190 191 194 211 212
+ 213 330 332 333 334 336 338 348 350 351
+ 352 354 356 366 368 369 370 372 374 505
+ 691 697 703 760 761 762 763
*.DEVICECLIMB
** N=789 EP=97 FDC=1597
X443 A3 gnd! B0 B2 B3 vdd! A2 A1 B1 50
+ A0 46 72 48 53 65 51 73 multiplier $T=1090 33260 0 0 $X=750 $Y=33040
X444 63 Cin vdd! gnd! A8 65 48 68 61 58
+ 56 49 54 55 73 51 72 57 53 50
+ 46 64 69 A9 59 67 47 52 66 71
+ 60 62 70 74 141 211 108 113 130 139
+ 140 158 159 176 185 190 191 194 212 213
+ 760 761 762 763 10badder $T=-50390 53780 1 0 $X=-110 $Y=0
X445 vdd! CLK gnd! RST A3 A_reg3 90 86 91 87
+ 506 88 508 84 85 89 92 ph1p3_MSDFF $T=1140 62320 0 0 $X=1140 $Y=58560
X446 vdd! CLK gnd! RST B0 B_reg0 81 77 82 78
+ 503 79 505 75 76 80 83 ph1p3_MSDFF $T=1140 69640 0 0 $X=1140 $Y=65880
X447 vdd! CLK gnd! RST A2 A_reg2 345 341 346 342
+ 692 343 694 339 340 344 347 ph1p3_MSDFF $T=11380 62320 0 0 $X=11380 $Y=58560
X448 vdd! CLK gnd! RST B1 B_reg1 336 332 337 333
+ 689 334 691 330 331 335 338 ph1p3_MSDFF $T=11380 69640 0 0 $X=11380 $Y=65880
X449 vdd! CLK gnd! RST A1 A_reg1 363 359 364 360
+ 698 361 700 357 358 362 365 ph1p3_MSDFF $T=21620 62320 0 0 $X=21620 $Y=58560
X450 vdd! CLK gnd! RST B2 B_reg2 354 350 355 351
+ 695 352 697 348 349 353 356 ph1p3_MSDFF $T=21620 69640 0 0 $X=21620 $Y=65880
X451 vdd! CLK gnd! RST A0 A_reg0 381 377 382 378
+ 704 379 706 375 376 380 383 ph1p3_MSDFF $T=31860 62320 0 0 $X=31860 $Y=58560
X452 vdd! CLK gnd! RST B3 B_reg3 372 368 373 369
+ 701 370 703 366 367 371 374 ph1p3_MSDFF $T=31860 69640 0 0 $X=31860 $Y=65880
X453 vdd! CLK gnd! RST 70 69 408 404 409 405
+ 713 406 715 402 403 407 410 ph1p3_MSDFF $T=37920 11080 0 0 $X=37920 $Y=7320
X454 vdd! CLK gnd! RST 64 63 399 395 400 396
+ 710 397 712 393 394 398 401 ph1p3_MSDFF $T=37920 18400 0 0 $X=37920 $Y=14640
X455 vdd! CLK gnd! RST 66 68 390 386 391 387
+ 707 388 709 384 385 389 392 ph1p3_MSDFF $T=37920 25720 0 0 $X=37920 $Y=21960
X456 vdd! CLK gnd! RST Sel Sel_reg 480 476 481 477
+ 737 478 739 474 475 479 482 ph1p3_MSDFF $T=48160 3760 0 0 $X=48160 $Y=0
X457 vdd! CLK gnd! RST 71 61 471 467 472 468
+ 734 469 736 465 466 470 473 ph1p3_MSDFF $T=48160 11080 0 0 $X=48160 $Y=7320
X458 vdd! CLK gnd! RST 60 58 462 458 463 459
+ 731 460 733 456 457 461 464 ph1p3_MSDFF $T=48160 18400 0 0 $X=48160 $Y=14640
X459 vdd! CLK gnd! RST 62 57 453 449 454 450
+ 728 451 730 447 448 452 455 ph1p3_MSDFF $T=48160 25720 0 0 $X=48160 $Y=21960
X460 vdd! CLK gnd! RST 67 56 444 440 445 441
+ 725 442 727 438 439 443 446 ph1p3_MSDFF $T=48160 33040 0 0 $X=48160 $Y=29280
X461 vdd! CLK gnd! RST 47 49 435 431 436 432
+ 722 433 724 429 430 434 437 ph1p3_MSDFF $T=48160 40360 0 0 $X=48160 $Y=36600
X462 vdd! CLK gnd! RST 52 54 426 422 427 423
+ 719 424 721 420 421 425 428 ph1p3_MSDFF $T=48160 47680 0 0 $X=48160 $Y=43920
X463 vdd! CLK gnd! RST 59 55 417 413 418 414
+ 716 415 718 411 412 416 419 ph1p3_MSDFF $T=48160 55000 0 0 $X=48160 $Y=51240
X465 Sel_reg 61 vdd! gnd! Sum_in6 Sum_out6 501 502 788 789 MUX_2to1___2X_ph2p2 $T=58160 11120 1 0 $X=58160 $Y=7320
X466 Sel_reg 69 vdd! gnd! Sum_in9 Sum_out9 499 500 786 787 MUX_2to1___2X_ph2p2 $T=58160 11080 0 0 $X=58160 $Y=11080
X467 Sel_reg 58 vdd! gnd! Sum_in5 Sum_out5 497 498 784 785 MUX_2to1___2X_ph2p2 $T=58160 18440 1 0 $X=58160 $Y=14640
X468 Sel_reg 63 vdd! gnd! Sum_in8 Sum_out8 495 496 782 783 MUX_2to1___2X_ph2p2 $T=58160 18400 0 0 $X=58160 $Y=18400
X469 Sel_reg 57 vdd! gnd! Sum_in4 Sum_out4 493 494 780 781 MUX_2to1___2X_ph2p2 $T=58160 25760 1 0 $X=58160 $Y=21960
X470 Sel_reg 68 vdd! gnd! Sum_in7 Sum_out7 491 492 778 779 MUX_2to1___2X_ph2p2 $T=58160 25720 0 0 $X=58160 $Y=25720
X471 Sel_reg 56 vdd! gnd! Sum_in3 Sum_out3 489 490 776 777 MUX_2to1___2X_ph2p2 $T=58160 33080 1 0 $X=58160 $Y=29280
X472 Sel_reg 49 vdd! gnd! Sum_in2 Sum_out2 487 488 774 775 MUX_2to1___2X_ph2p2 $T=58160 40400 1 0 $X=58160 $Y=36600
X473 Sel_reg 54 vdd! gnd! Sum_in1 Sum_out1 485 486 772 773 MUX_2to1___2X_ph2p2 $T=58160 47720 1 0 $X=58160 $Y=43920
X474 Sel_reg 55 vdd! gnd! Sum_in0 Sum_out0 483 484 770 771 MUX_2to1___2X_ph2p2 $T=58160 55040 1 0 $X=58160 $Y=51240
M0 87 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=59450 $dt=1
M1 90 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=64750 $dt=1
M2 78 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=66770 $dt=1
M3 84 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3250 $Y=64780 $dt=1
M4 85 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=59420 $dt=1
M5 76 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=66740 $dt=1
M6 86 CLK A3 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4430 $Y=64780 $dt=1
M7 91 CLK 506 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=59660 $dt=1
M8 82 CLK 503 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=66980 $dt=1
M9 88 86 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5630 $Y=64690 $dt=1
M10 506 A_reg3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=59450 $dt=1
M11 503 B_reg0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=66770 $dt=1
M12 88 87 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6870 $Y=64700 $dt=1
M13 89 90 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=59420 $dt=1
M14 80 81 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=66740 $dt=1
M15 508 88 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8120 $Y=64750 $dt=1
M16 91 90 88 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=59660 $dt=1
M17 82 81 79 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=66980 $dt=1
M18 92 90 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9450 $Y=64780 $dt=1
M19 A_reg3 91 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=59450 $dt=1
M20 B_reg0 82 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=66770 $dt=1
M21 86 90 508 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=10630 $Y=64780 $dt=1
M22 342 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=59450 $dt=1
M23 345 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=64750 $dt=1
M24 333 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=66770 $dt=1
M25 339 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13490 $Y=64780 $dt=1
M26 340 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=59420 $dt=1
M27 331 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=66740 $dt=1
M28 341 CLK A2 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=14670 $Y=64780 $dt=1
M29 346 CLK 692 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=59660 $dt=1
M30 337 CLK 689 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=66980 $dt=1
M31 343 341 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=15870 $Y=64690 $dt=1
M32 692 A_reg2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=59450 $dt=1
M33 689 B_reg1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=66770 $dt=1
M34 343 342 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17110 $Y=64700 $dt=1
M35 344 345 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=59420 $dt=1
M36 335 336 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=66740 $dt=1
M37 694 343 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18360 $Y=64750 $dt=1
M38 346 345 343 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=59660 $dt=1
M39 337 336 334 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=66980 $dt=1
M40 347 345 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=19690 $Y=64780 $dt=1
M41 A_reg2 346 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=59450 $dt=1
M42 B_reg1 337 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=66770 $dt=1
M43 341 345 694 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=20870 $Y=64780 $dt=1
M44 360 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=59450 $dt=1
M45 363 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=64750 $dt=1
M46 351 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=66770 $dt=1
M47 357 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=23730 $Y=64780 $dt=1
M48 358 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=59420 $dt=1
M49 349 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=66740 $dt=1
M50 359 CLK A1 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=24910 $Y=64780 $dt=1
M51 364 CLK 698 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=59660 $dt=1
M52 355 CLK 695 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=66980 $dt=1
M53 361 359 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26110 $Y=64690 $dt=1
M54 698 A_reg1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=59450 $dt=1
M55 695 B_reg2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=66770 $dt=1
M56 361 360 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27350 $Y=64700 $dt=1
M57 362 363 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=59420 $dt=1
M58 353 354 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=66740 $dt=1
M59 700 361 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28600 $Y=64750 $dt=1
M60 364 363 361 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=59660 $dt=1
M61 355 354 352 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=66980 $dt=1
M62 365 363 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=29930 $Y=64780 $dt=1
M63 A_reg1 364 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=59450 $dt=1
M64 B_reg2 355 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=66770 $dt=1
M65 359 363 700 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31110 $Y=64780 $dt=1
M66 378 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=59450 $dt=1
M67 381 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=64750 $dt=1
M68 369 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=66770 $dt=1
M69 375 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=33970 $Y=64780 $dt=1
M70 376 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=59420 $dt=1
M71 367 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=66740 $dt=1
M72 377 CLK A0 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35150 $Y=64780 $dt=1
M73 382 CLK 704 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=59660 $dt=1
M74 373 CLK 701 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=66980 $dt=1
M75 379 377 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36350 $Y=64690 $dt=1
M76 704 A_reg0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=37440 $Y=59450 $dt=1
M77 701 B_reg3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=37440 $Y=66770 $dt=1
M78 379 378 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37590 $Y=64700 $dt=1
M79 405 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=8210 $dt=1
M80 408 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=13510 $dt=1
M81 396 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=15530 $dt=1
M82 399 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=20830 $dt=1
M83 387 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=22850 $dt=1
M84 390 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=28150 $dt=1
M85 380 381 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=38770 $Y=59420 $dt=1
M86 371 372 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=38770 $Y=66740 $dt=1
M87 706 379 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=38840 $Y=64750 $dt=1
M88 382 381 379 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=39950 $Y=59660 $dt=1
M89 373 372 370 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=39950 $Y=66980 $dt=1
M90 402 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=13540 $dt=1
M91 393 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=20860 $dt=1
M92 384 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=40030 $Y=28180 $dt=1
M93 383 381 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40170 $Y=64780 $dt=1
M94 403 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=41030 $Y=8180 $dt=1
M95 394 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=15500 $dt=1
M96 385 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=22820 $dt=1
M97 404 CLK 70 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=13540 $dt=1
M98 395 CLK 64 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=20860 $dt=1
M99 386 CLK 66 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=41210 $Y=28180 $dt=1
M100 A_reg0 382 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=41240 $Y=59450 $dt=1
M101 B_reg3 373 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=41240 $Y=66770 $dt=1
M102 377 381 706 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41350 $Y=64780 $dt=1
M103 409 CLK 713 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=42210 $Y=8420 $dt=1
M104 400 CLK 710 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=15740 $dt=1
M105 391 CLK 707 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=23060 $dt=1
M106 406 404 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=13450 $dt=1
M107 397 395 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=20770 $dt=1
M108 388 386 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42410 $Y=28090 $dt=1
M109 713 69 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=43500 $Y=8210 $dt=1
M110 710 63 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=15530 $dt=1
M111 707 68 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=22850 $dt=1
M112 406 405 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=13460 $dt=1
M113 397 396 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=20780 $dt=1
M114 388 387 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43650 $Y=28100 $dt=1
M115 407 408 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=44830 $Y=8180 $dt=1
M116 398 399 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=15500 $dt=1
M117 389 390 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=22820 $dt=1
M118 715 406 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=13510 $dt=1
M119 712 397 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=20830 $dt=1
M120 709 388 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=44900 $Y=28150 $dt=1
M121 409 408 406 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=46010 $Y=8420 $dt=1
M122 400 399 397 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=15740 $dt=1
M123 391 390 388 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=23060 $dt=1
M124 410 408 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=13540 $dt=1
M125 401 399 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=20860 $dt=1
M126 392 390 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=46230 $Y=28180 $dt=1
M127 69 409 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=47300 $Y=8210 $dt=1
M128 63 400 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=15530 $dt=1
M129 68 391 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=22850 $dt=1
M130 404 408 715 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=13540 $dt=1
M131 395 399 712 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=20860 $dt=1
M132 386 390 709 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=47410 $Y=28180 $dt=1
M133 477 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=890 $dt=1
M134 480 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=6190 $dt=1
M135 468 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=8210 $dt=1
M136 471 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=13510 $dt=1
M137 459 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=15530 $dt=1
M138 462 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=20830 $dt=1
M139 450 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=22850 $dt=1
M140 453 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=28150 $dt=1
M141 441 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=30170 $dt=1
M142 444 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=35470 $dt=1
M143 432 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=37490 $dt=1
M144 435 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=42790 $dt=1
M145 423 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=44810 $dt=1
M146 426 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=50110 $dt=1
M147 414 RST vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=52130 $dt=1
M148 417 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=57430 $dt=1
M149 474 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=6220 $dt=1
M150 465 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=13540 $dt=1
M151 456 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=20860 $dt=1
M152 447 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=28180 $dt=1
M153 438 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=35500 $dt=1
M154 429 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=42820 $dt=1
M155 420 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=50140 $dt=1
M156 411 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=50270 $Y=57460 $dt=1
M157 475 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=51270 $Y=860 $dt=1
M158 466 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=8180 $dt=1
M159 457 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=15500 $dt=1
M160 448 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=22820 $dt=1
M161 439 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=30140 $dt=1
M162 430 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=37460 $dt=1
M163 421 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=44780 $dt=1
M164 412 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=52100 $dt=1
M165 476 CLK Sel vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=6220 $dt=1
M166 467 CLK 71 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=13540 $dt=1
M167 458 CLK 60 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=20860 $dt=1
M168 449 CLK 62 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=28180 $dt=1
M169 440 CLK 67 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=35500 $dt=1
M170 431 CLK 47 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=42820 $dt=1
M171 422 CLK 52 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=50140 $dt=1
M172 413 CLK 59 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=51450 $Y=57460 $dt=1
M173 481 CLK 737 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=52450 $Y=1100 $dt=1
M174 472 CLK 734 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=8420 $dt=1
M175 463 CLK 731 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=15740 $dt=1
M176 454 CLK 728 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=23060 $dt=1
M177 445 CLK 725 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=30380 $dt=1
M178 436 CLK 722 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=37700 $dt=1
M179 427 CLK 719 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=45020 $dt=1
M180 418 CLK 716 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=52340 $dt=1
M181 478 476 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=6130 $dt=1
M182 469 467 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=13450 $dt=1
M183 460 458 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=20770 $dt=1
M184 451 449 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=28090 $dt=1
M185 442 440 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=35410 $dt=1
M186 433 431 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=42730 $dt=1
M187 424 422 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=50050 $dt=1
M188 415 413 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=52650 $Y=57370 $dt=1
M189 737 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=53740 $Y=890 $dt=1
M190 734 61 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=8210 $dt=1
M191 731 58 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=15530 $dt=1
M192 728 57 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=22850 $dt=1
M193 725 56 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=30170 $dt=1
M194 722 49 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=37490 $dt=1
M195 719 54 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=44810 $dt=1
M196 716 55 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=52130 $dt=1
M197 478 477 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=6140 $dt=1
M198 469 468 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=13460 $dt=1
M199 460 459 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=20780 $dt=1
M200 451 450 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=28100 $dt=1
M201 442 441 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=35420 $dt=1
M202 433 432 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=42740 $dt=1
M203 424 423 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=50060 $dt=1
M204 415 414 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=53890 $Y=57380 $dt=1
M205 479 480 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=55070 $Y=860 $dt=1
M206 470 471 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=8180 $dt=1
M207 461 462 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=15500 $dt=1
M208 452 453 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=22820 $dt=1
M209 443 444 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=30140 $dt=1
M210 434 435 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=37460 $dt=1
M211 425 426 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=44780 $dt=1
M212 416 417 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=52100 $dt=1
M213 739 478 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=6190 $dt=1
M214 736 469 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=13510 $dt=1
M215 733 460 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=20830 $dt=1
M216 730 451 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=28150 $dt=1
M217 727 442 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=35470 $dt=1
M218 724 433 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=42790 $dt=1
M219 721 424 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=50110 $dt=1
M220 718 415 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=55140 $Y=57430 $dt=1
M221 481 480 478 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=56250 $Y=1100 $dt=1
M222 472 471 469 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=8420 $dt=1
M223 463 462 460 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=15740 $dt=1
M224 454 453 451 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=23060 $dt=1
M225 445 444 442 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=30380 $dt=1
M226 436 435 433 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=37700 $dt=1
M227 427 426 424 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=45020 $dt=1
M228 418 417 415 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=52340 $dt=1
M229 482 480 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=6220 $dt=1
M230 473 471 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=13540 $dt=1
M231 464 462 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=20860 $dt=1
M232 455 453 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=28180 $dt=1
M233 446 444 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=35500 $dt=1
M234 437 435 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=42820 $dt=1
M235 428 426 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=50140 $dt=1
M236 419 417 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=56470 $Y=57460 $dt=1
M237 Sel_reg 481 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=57540 $Y=890 $dt=1
M238 61 472 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=8210 $dt=1
M239 58 463 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=15530 $dt=1
M240 57 454 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=22850 $dt=1
M241 56 445 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=30170 $dt=1
M242 49 436 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=37490 $dt=1
M243 54 427 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=44810 $dt=1
M244 55 418 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=52130 $dt=1
M245 476 480 739 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=6220 $dt=1
M246 467 471 736 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=13540 $dt=1
M247 458 462 733 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=20860 $dt=1
M248 449 453 730 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=28180 $dt=1
M249 440 444 727 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=35500 $dt=1
M250 431 435 724 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=42820 $dt=1
M251 422 426 721 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=50140 $dt=1
M252 413 417 718 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=57650 $Y=57460 $dt=1
M253 501 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=8270 $dt=1
M254 499 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=13450 $dt=1
M255 497 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=15590 $dt=1
M256 495 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=20770 $dt=1
M257 493 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=22910 $dt=1
M258 491 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=28090 $dt=1
M259 489 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=30230 $dt=1
M260 487 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=37550 $dt=1
M261 485 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=44870 $dt=1
M262 483 Sel_reg vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=52190 $dt=1
M263 788 61 502 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=8060 $dt=1
M264 786 69 500 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=13180 $dt=1
M265 784 58 498 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=15380 $dt=1
M266 782 63 496 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=20500 $dt=1
M267 780 57 494 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=22700 $dt=1
M268 778 68 492 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=27820 $dt=1
M269 776 56 490 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=30020 $dt=1
M270 774 49 488 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=37340 $dt=1
M271 772 54 486 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=44660 $dt=1
M272 770 55 484 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=51980 $dt=1
M273 vdd! Sel_reg 788 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=8060 $dt=1
M274 vdd! Sel_reg 786 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=13180 $dt=1
M275 vdd! Sel_reg 784 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=15380 $dt=1
M276 vdd! Sel_reg 782 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=20500 $dt=1
M277 vdd! Sel_reg 780 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=22700 $dt=1
M278 vdd! Sel_reg 778 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=27820 $dt=1
M279 vdd! Sel_reg 776 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=30020 $dt=1
M280 vdd! Sel_reg 774 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=37340 $dt=1
M281 vdd! Sel_reg 772 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=44660 $dt=1
M282 vdd! Sel_reg 770 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=51980 $dt=1
M283 789 501 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=8130 $dt=1
M284 787 499 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=13110 $dt=1
M285 785 497 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=15450 $dt=1
M286 783 495 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=20430 $dt=1
M287 781 493 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=22770 $dt=1
M288 779 491 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=27750 $dt=1
M289 777 489 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=30090 $dt=1
M290 775 487 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=37410 $dt=1
M291 773 485 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=44730 $dt=1
M292 771 483 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=52050 $dt=1
M293 502 Sum_in6 789 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=8130 $dt=1
M294 500 Sum_in9 787 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=13110 $dt=1
M295 498 Sum_in5 785 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=15450 $dt=1
M296 496 Sum_in8 783 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=20430 $dt=1
M297 494 Sum_in4 781 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=22770 $dt=1
M298 492 Sum_in7 779 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=27750 $dt=1
M299 490 Sum_in3 777 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=30090 $dt=1
M300 488 Sum_in2 775 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=37410 $dt=1
M301 486 Sum_in1 773 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=44730 $dt=1
M302 484 Sum_in0 771 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=52050 $dt=1
M303 Sum_out6 502 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=8120 $dt=1
M304 Sum_out9 500 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=13120 $dt=1
M305 Sum_out5 498 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=15440 $dt=1
M306 Sum_out8 496 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=20440 $dt=1
M307 Sum_out4 494 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=22760 $dt=1
M308 Sum_out7 492 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=27760 $dt=1
M309 Sum_out3 490 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=30080 $dt=1
M310 Sum_out2 488 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=37400 $dt=1
M311 Sum_out1 486 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=44720 $dt=1
M312 Sum_out0 484 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=52040 $dt=1
.ends ph2p2_processing_element

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p3_Matrix_vector_Multiplication              *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p3_Matrix_vector_Multiplication A3_3 A2_3 A1_3 A0_3 B_reg0 A3_1 gnd! A3_reg3 Cin3 CLK
+ RST A3_8 vdd! A2_1 A2_reg3 Cin2 A2_8 A1_1 A1_reg3 Cin1
+ A1_8 A0_1 B0_1 A0_reg3 B0_0 B0_2 B0_3 Cin0 A0_8 A3_2
+ A2_2 A1_2 A0_2 B_reg1 A3_reg2 A3_0 A2_reg2 A2_0 A1_reg2 A1_0
+ A0_reg2 A0_0 B_reg2 A0_reg1 A1_reg1 A2_reg1 A3_reg1 A3_9 A2_9 A1_9
+ A0_9 B_reg3 A3_reg0 A2_reg0 A1_reg0 A0_reg0 Sel3 Sel2 Sel1 Sel0
+ Sel0_reg Sel1_reg Sel2_reg Sel3_reg Sum_in0 Sum_in1 Sum_in2 Sum_in3 Sum_in7 Sum_in4
+ Sum_in8 Sum_in5 Sum_in9 Sum_in6 Sum_out0 Sum_out2 Sum_out9 Sum_out1 Sum_out3 Sum_out7
+ Sum_out4 Sum_out8 Sum_out5 Sum_out6
** N=2678 EP=84 FDC=6648
X324 A3_3 115 124 121 gnd! RST CLK Cin3 A3_8 vdd!
+ 118 A3_reg3 B_reg0 A3_1 A3_2 A3_0 B_reg1 A3_reg2 A3_9 B_reg2
+ A3_reg1 A3_reg0 B_reg3 Sel3 Sel3_reg 100 106 85 97 112
+ 101 88 109 94 91 Sum_in6 Sum_in9 Sum_in5 Sum_in8 Sum_in4
+ Sum_in7 Sum_in3 Sum_in2 Sum_in1 Sum_in0 1232 2362 1377 2466 2663
+ 2599 2600 2601 2602 2666 1244 1256 1291 1302 1306
+ 1316 1353 1354 1397 1402 1420 1425 1431 1459 1477
+ 1478 2668 2603 2604 2605 2606 2670 2671 2607 2608
+ 2609 2610 2674 2676 2611 2612 2613 2614 2678 2665
+ 2669 2673 2677 2664 2667 2672 2675 ph2p2_processing_element $T=370 -60 0 0 $X=260 $Y=-60
X325 A2_3 116 125 122 gnd! RST CLK Cin2 A2_8 vdd!
+ 119 A2_reg3 115 A2_1 A2_2 A2_0 118 A2_reg2 A2_9 124
+ A2_reg1 A2_reg0 121 Sel2 Sel2_reg 102 107 86 98 113
+ 103 89 110 95 92 94 97 100 101 88
+ 91 85 109 112 106 867 2121 1012 2225 2647
+ 2583 2584 2585 2586 2650 879 891 926 937 941
+ 951 988 989 1032 1037 1055 1060 1066 1094 1112
+ 1113 2652 2587 2588 2589 2590 2654 2655 2591 2592
+ 2593 2594 2658 2660 2595 2596 2597 2598 2662 2649
+ 2653 2657 2661 2648 2651 2656 2659 ph2p2_processing_element $T=370 73140 0 0 $X=260 $Y=73140
X326 A1_3 117 126 123 gnd! RST CLK Cin1 A1_8 vdd!
+ 120 A1_reg3 116 A1_1 A1_2 A1_0 119 A1_reg2 A1_9 125
+ A1_reg1 A1_reg0 122 Sel1 Sel1_reg 104 108 87 99 114
+ 105 90 111 96 93 95 98 102 103 89
+ 92 86 110 113 107 502 1880 647 1984 2631
+ 2567 2568 2569 2570 2634 514 526 561 572 576
+ 586 623 624 667 672 690 695 701 729 747
+ 748 2636 2571 2572 2573 2574 2638 2639 2575 2576
+ 2577 2578 2642 2644 2579 2580 2581 2582 2646 2633
+ 2637 2641 2645 2632 2635 2640 2643 ph2p2_processing_element $T=370 146340 0 0 $X=260 $Y=146340
X327 A0_3 B0_0 B0_2 B0_3 gnd! RST CLK Cin0 A0_8 vdd!
+ B0_1 A0_reg3 117 A0_1 A0_2 A0_0 120 A0_reg2 A0_9 126
+ A0_reg1 A0_reg0 123 Sel0 Sel0_reg Sum_out5 Sum_out0 Sum_out3 Sum_out9 Sum_out1
+ Sum_out8 Sum_out4 Sum_out2 Sum_out6 Sum_out7 96 99 104 105 90
+ 93 87 111 114 108 137 1639 282 1743 2615
+ 2551 2552 2553 2554 2618 149 161 196 207 211
+ 221 258 259 302 307 325 330 336 364 382
+ 383 2620 2555 2556 2557 2558 2622 2623 2559 2560
+ 2561 2562 2626 2628 2563 2564 2565 2566 2630 2617
+ 2621 2625 2629 2616 2619 2624 2627 ph2p2_processing_element $T=370 219540 0 0 $X=260 $Y=219540
M0 2602 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=72010 $dt=1
M1 2586 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=145210 $dt=1
M2 2570 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=218410 $dt=1
M3 2554 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=2290 $Y=291610 $dt=1
M4 1256 1232 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.8911 scb=0.00996238 scc=0.000256798 $X=2380 $Y=920 $dt=1
M5 891 867 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=74120 $dt=1
M6 526 502 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=147320 $dt=1
M7 161 137 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=220520 $dt=1
M8 2663 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=72040 $dt=1
M9 2647 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=145240 $dt=1
M10 2631 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=218440 $dt=1
M11 2615 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=3620 $Y=291640 $dt=1
M12 2664 1232 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=3710 $Y=680 $dt=1
M13 2648 867 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=73880 $dt=1
M14 2632 502 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=147080 $dt=1
M15 2616 137 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=220280 $dt=1
M16 1291 1244 2664 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=4680 $Y=620 $dt=1
M17 926 879 2648 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=73820 $dt=1
M18 561 514 2632 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=147020 $dt=1
M19 196 149 2616 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=220220 $dt=1
M20 2599 CLK 115 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=72040 $dt=1
M21 2583 CLK 116 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=145240 $dt=1
M22 2567 CLK 117 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=218440 $dt=1
M23 2551 CLK B0_0 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=4800 $Y=291640 $dt=1
M24 1291 1256 2664 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=5640 $Y=620 $dt=1
M25 926 891 2648 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=73820 $dt=1
M26 561 526 2632 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=147020 $dt=1
M27 196 161 2616 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=220220 $dt=1
M28 2601 2599 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=71950 $dt=1
M29 2585 2583 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=145150 $dt=1
M30 2569 2567 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=218350 $dt=1
M31 2553 2551 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=6000 $Y=291550 $dt=1
M32 2664 A3_8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=6600 $Y=620 $dt=1
M33 2648 A2_8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=73820 $dt=1
M34 2632 A1_8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=147020 $dt=1
M35 2616 A0_8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=220220 $dt=1
M36 2601 2600 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=71960 $dt=1
M37 2585 2584 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=145160 $dt=1
M38 2569 2568 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=218360 $dt=1
M39 2553 2552 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=7240 $Y=291560 $dt=1
M40 1302 1316 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=8260 $Y=920 $dt=1
M41 937 951 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=74120 $dt=1
M42 572 586 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=147320 $dt=1
M43 207 221 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=220520 $dt=1
M44 2665 2601 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=72010 $dt=1
M45 2649 2585 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=145210 $dt=1
M46 2633 2569 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=218410 $dt=1
M47 2617 2553 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=8490 $Y=291610 $dt=1
M48 1306 1291 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=9220 $Y=920 $dt=1
M49 941 926 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=74120 $dt=1
M50 576 561 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=147320 $dt=1
M51 211 196 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=220520 $dt=1
M52 2666 2602 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=72040 $dt=1
M53 2650 2586 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=145240 $dt=1
M54 2634 2570 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=218440 $dt=1
M55 2618 2554 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=9820 $Y=291640 $dt=1
M56 2667 1291 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=10550 $Y=680 $dt=1
M57 2651 926 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=73880 $dt=1
M58 2635 561 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=147080 $dt=1
M59 2619 196 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=220280 $dt=1
M60 2599 2602 2665 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=72040 $dt=1
M61 2583 2586 2649 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=145240 $dt=1
M62 2567 2570 2633 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=218440 $dt=1
M63 2551 2554 2617 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=11000 $Y=291640 $dt=1
M64 2362 1302 2667 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=11520 $Y=620 $dt=1
M65 2121 937 2651 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=73820 $dt=1
M66 1880 572 2635 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=147020 $dt=1
M67 1639 207 2619 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=220220 $dt=1
M68 2362 1306 2667 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=12480 $Y=620 $dt=1
M69 2121 941 2651 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=73820 $dt=1
M70 1880 576 2635 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=147020 $dt=1
M71 1639 211 2619 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=220220 $dt=1
M72 2606 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=72010 $dt=1
M73 2590 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=145210 $dt=1
M74 2574 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=218410 $dt=1
M75 2558 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=12530 $Y=291610 $dt=1
M76 2667 1316 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=13440 $Y=620 $dt=1
M77 2651 951 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=73820 $dt=1
M78 2635 586 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=147020 $dt=1
M79 2619 221 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=220220 $dt=1
M80 2668 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=72040 $dt=1
M81 2652 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=145240 $dt=1
M82 2636 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=218440 $dt=1
M83 2620 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=13860 $Y=291640 $dt=1
M84 2603 CLK 118 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=72040 $dt=1
M85 2587 CLK 119 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=145240 $dt=1
M86 2571 CLK 120 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=218440 $dt=1
M87 2555 CLK B0_1 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=15040 $Y=291640 $dt=1
M88 1353 1316 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=15510 $Y=650 $dt=1
M89 988 951 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=73850 $dt=1
M90 623 586 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=147050 $dt=1
M91 258 221 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=220250 $dt=1
M92 vdd! 1291 1353 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=15920 $Y=650 $dt=1
M93 vdd! 926 988 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=73850 $dt=1
M94 vdd! 561 623 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=147050 $dt=1
M95 vdd! 196 258 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=220250 $dt=1
M96 2605 2603 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=71950 $dt=1
M97 2589 2587 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=145150 $dt=1
M98 2573 2571 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=218350 $dt=1
M99 2557 2555 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=16240 $Y=291550 $dt=1
M100 2605 2604 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=71960 $dt=1
M101 2589 2588 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=145160 $dt=1
M102 2573 2572 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=218360 $dt=1
M103 2557 2556 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=17480 $Y=291560 $dt=1
M104 1354 A3_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=18490 $Y=910 $dt=1
M105 989 A2_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=74110 $dt=1
M106 624 A1_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=147310 $dt=1
M107 259 A0_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=220510 $dt=1
M108 2669 2605 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=72010 $dt=1
M109 2653 2589 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=145210 $dt=1
M110 2637 2573 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=218410 $dt=1
M111 2621 2557 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=18730 $Y=291610 $dt=1
M112 vdd! 1232 1354 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=18900 $Y=910 $dt=1
M113 vdd! 867 989 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=74110 $dt=1
M114 vdd! 502 624 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=147310 $dt=1
M115 vdd! 137 259 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=220510 $dt=1
M116 2670 2606 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=72040 $dt=1
M117 2654 2590 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=145240 $dt=1
M118 2638 2574 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=218440 $dt=1
M119 2622 2558 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=20060 $Y=291640 $dt=1
M120 2603 2606 2669 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=72040 $dt=1
M121 2587 2590 2653 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=145240 $dt=1
M122 2571 2574 2637 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=218440 $dt=1
M123 2555 2558 2621 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=21240 $Y=291640 $dt=1
M124 1459 1353 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=21330 $Y=910 $dt=1
M125 1094 988 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=74110 $dt=1
M126 729 623 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=147310 $dt=1
M127 364 258 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=220510 $dt=1
M128 vdd! 1354 1459 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=21740 $Y=910 $dt=1
M129 vdd! 989 1094 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=74110 $dt=1
M130 vdd! 624 729 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=147310 $dt=1
M131 vdd! 259 364 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=220510 $dt=1
M132 2610 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=72010 $dt=1
M133 2594 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=145210 $dt=1
M134 2578 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=218410 $dt=1
M135 2562 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=22770 $Y=291610 $dt=1
M136 1397 A3_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=23380 $Y=920 $dt=1
M137 1032 A2_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=74120 $dt=1
M138 667 A1_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=147320 $dt=1
M139 302 A0_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=220520 $dt=1
M140 2671 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=72040 $dt=1
M141 2655 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=145240 $dt=1
M142 2639 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=218440 $dt=1
M143 2623 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=24100 $Y=291640 $dt=1
M144 1402 1377 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=24340 $Y=920 $dt=1
M145 1037 1012 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=74120 $dt=1
M146 672 647 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=147320 $dt=1
M147 307 282 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=220520 $dt=1
M148 2607 CLK 124 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=72040 $dt=1
M149 2591 CLK 125 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=145240 $dt=1
M150 2575 CLK 126 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=218440 $dt=1
M151 2559 CLK B0_2 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=25280 $Y=291640 $dt=1
M152 2672 1377 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=25670 $Y=680 $dt=1
M153 2656 1012 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=73880 $dt=1
M154 2640 647 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=147080 $dt=1
M155 2624 282 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=220280 $dt=1
M156 2609 2607 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=71950 $dt=1
M157 2593 2591 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=145150 $dt=1
M158 2577 2575 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=218350 $dt=1
M159 2561 2559 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=26480 $Y=291550 $dt=1
M160 1420 1397 2672 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=26640 $Y=620 $dt=1
M161 1055 1032 2656 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=73820 $dt=1
M162 690 667 2640 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=147020 $dt=1
M163 325 302 2624 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=220220 $dt=1
M164 1420 1402 2672 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=27600 $Y=620 $dt=1
M165 1055 1037 2656 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=73820 $dt=1
M166 690 672 2640 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=147020 $dt=1
M167 325 307 2624 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=220220 $dt=1
M168 2609 2608 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=71960 $dt=1
M169 2593 2592 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=145160 $dt=1
M170 2577 2576 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=218360 $dt=1
M171 2561 2560 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=27720 $Y=291560 $dt=1
M172 2672 A3_9 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=28560 $Y=620 $dt=1
M173 2656 A2_9 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=73820 $dt=1
M174 2640 A1_9 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=147020 $dt=1
M175 2624 A0_9 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=220220 $dt=1
M176 2673 2609 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=72010 $dt=1
M177 2657 2593 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=145210 $dt=1
M178 2641 2577 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=218410 $dt=1
M179 2625 2561 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=28970 $Y=291610 $dt=1
M180 1425 1459 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=30220 $Y=920 $dt=1
M181 1060 1094 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=74120 $dt=1
M182 695 729 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=147320 $dt=1
M183 330 364 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=220520 $dt=1
M184 2674 2610 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=72040 $dt=1
M185 2658 2594 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=145240 $dt=1
M186 2642 2578 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=218440 $dt=1
M187 2626 2562 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=30300 $Y=291640 $dt=1
M188 1431 1420 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=31180 $Y=920 $dt=1
M189 1066 1055 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=74120 $dt=1
M190 701 690 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=147320 $dt=1
M191 336 325 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=220520 $dt=1
M192 2607 2610 2673 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=72040 $dt=1
M193 2591 2594 2657 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=145240 $dt=1
M194 2575 2578 2641 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=218440 $dt=1
M195 2559 2562 2625 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=31480 $Y=291640 $dt=1
M196 2675 1420 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=32510 $Y=680 $dt=1
M197 2659 1055 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=73880 $dt=1
M198 2643 690 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=147080 $dt=1
M199 2627 325 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=220280 $dt=1
M200 2614 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=72010 $dt=1
M201 2598 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=145210 $dt=1
M202 2582 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=218410 $dt=1
M203 2566 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=33010 $Y=291610 $dt=1
M204 2466 1425 2675 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=33480 $Y=620 $dt=1
M205 2225 1060 2659 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=73820 $dt=1
M206 1984 695 2643 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=147020 $dt=1
M207 1743 330 2627 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=220220 $dt=1
M208 2676 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=72040 $dt=1
M209 2660 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=145240 $dt=1
M210 2644 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=218440 $dt=1
M211 2628 CLK vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=34340 $Y=291640 $dt=1
M212 2466 1431 2675 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=34440 $Y=620 $dt=1
M213 2225 1066 2659 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=73820 $dt=1
M214 1984 701 2643 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=147020 $dt=1
M215 1743 336 2627 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=220220 $dt=1
M216 2675 1459 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=35400 $Y=620 $dt=1
M217 2659 1094 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=73820 $dt=1
M218 2643 729 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=147020 $dt=1
M219 2627 364 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=220220 $dt=1
M220 2611 CLK 121 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=72040 $dt=1
M221 2595 CLK 122 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=145240 $dt=1
M222 2579 CLK 123 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=218440 $dt=1
M223 2563 CLK B0_3 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=35520 $Y=291640 $dt=1
M224 2613 2611 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=71950 $dt=1
M225 2597 2595 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=145150 $dt=1
M226 2581 2579 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=218350 $dt=1
M227 2565 2563 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=36720 $Y=291550 $dt=1
M228 1477 1459 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=37470 $Y=650 $dt=1
M229 1112 1094 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=73850 $dt=1
M230 747 729 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=147050 $dt=1
M231 382 364 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=220250 $dt=1
M232 vdd! 1420 1477 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=37880 $Y=650 $dt=1
M233 vdd! 1055 1112 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=73850 $dt=1
M234 vdd! 690 747 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=147050 $dt=1
M235 vdd! 325 382 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=220250 $dt=1
M236 2613 2612 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=71960 $dt=1
M237 2597 2596 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=145160 $dt=1
M238 2581 2580 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=218360 $dt=1
M239 2565 2564 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=37960 $Y=291560 $dt=1
M240 2677 2613 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=72010 $dt=1
M241 2661 2597 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=145210 $dt=1
M242 2645 2581 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=218410 $dt=1
M243 2629 2565 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=39210 $Y=291610 $dt=1
M244 1478 A3_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=40450 $Y=910 $dt=1
M245 1113 A2_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=74110 $dt=1
M246 748 A1_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=147310 $dt=1
M247 383 A0_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=220510 $dt=1
M248 2678 2614 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=72040 $dt=1
M249 2662 2598 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=145240 $dt=1
M250 2646 2582 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=218440 $dt=1
M251 2630 2566 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=40540 $Y=291640 $dt=1
M252 vdd! 1377 1478 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=40860 $Y=910 $dt=1
M253 vdd! 1012 1113 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=74110 $dt=1
M254 vdd! 647 748 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=147310 $dt=1
M255 vdd! 282 383 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=220510 $dt=1
M256 2611 2614 2677 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=72040 $dt=1
M257 2595 2598 2661 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=145240 $dt=1
M258 2579 2582 2645 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=218440 $dt=1
M259 2563 2566 2629 vdd! g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=41720 $Y=291640 $dt=1
.ends ph2p3_Matrix_vector_Multiplication

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph3_sytolic_array                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph3_sytolic_array A0_0 A0_0_8 A0_0_9 A0_1 A0_1_8 A0_1_9 A0_2 A0_2_8 A0_2_9 A0_3
+ A0_3_8 A0_3_9 A0_reg0 A0_reg1 A0_reg2 A0_reg3 A1_0 A1_0_8 A1_0_9 A1_1
+ A1_1_8 A1_1_9 A1_2 A1_2_8 A1_2_9 A1_3 A1_3_8 A1_3_9 A1_reg0 A1_reg1
+ A1_reg2 A1_reg3 A2_0 A2_0_8 A2_0_9 A2_1 A2_1_8 A2_1_9 A2_2 A2_2_8
+ A2_2_9 A2_3 A2_3_8 A2_3_9 A2_reg0 A2_reg1 A2_reg2 A2_reg3 A3_0 A3_0_8
+ A3_0_9 A3_1 A3_1_8 A3_1_9 A3_2 A3_2_8 A3_2_9 A3_3 A3_3_8 A3_3_9
+ A3_reg0 A3_reg1 A3_reg2 A3_reg3 B0_0 B0_1 B0_2 B0_3 B0_reg0 B0_reg1
+ B0_reg2 B0_reg3 B1_0 B1_1 B1_2 B1_3 B1_reg0 B1_reg1 B1_reg2 B1_reg3
+ B2_0 B2_1 B2_2 B2_3 B2_reg0 B2_reg1 B2_reg2 B2_reg3 B3_0 B3_1
+ B3_2 B3_3 B3_reg0 B3_reg1 B3_reg2 B3_reg3 CLK Cin0_0 Cin0_1 Cin0_2
+ Cin0_3 Cin1_0 Cin1_1 Cin1_2 Cin1_3 Cin2_0 Cin2_1 Cin2_2 Cin2_3 Cin3_0
+ Cin3_1 Cin3_2 Cin3_3 RST Sel0 Sel1 Sel2 Sel3 Sum0_in0 Sum0_in1
+ Sum0_in2 Sum0_in3 Sum0_in4 Sum0_in5 Sum0_in6 Sum0_in7 Sum0_in8 Sum0_in9 Sum0_out0 Sum0_out1
+ Sum0_out2 Sum0_out3 Sum0_out4 Sum0_out5 Sum0_out6 Sum0_out7 Sum0_out8 Sum0_out9 Sum1_in0 Sum1_in1
+ Sum1_in2 Sum1_in3 Sum1_in4 Sum1_in5 Sum1_in6 Sum1_in7 Sum1_in8 Sum1_in9 Sum1_out0 Sum1_out1
+ Sum1_out2 Sum1_out3 Sum1_out4 Sum1_out5 Sum1_out6 Sum1_out7 Sum1_out8 Sum1_out9 Sum2_in0 Sum2_in1
+ Sum2_in2 Sum2_in3 Sum2_in4 Sum2_in5 Sum2_in6 Sum2_in7 Sum2_in8 Sum2_in9 Sum2_out0 Sum2_out1
+ Sum2_out2 Sum2_out3 Sum2_out4 Sum2_out5 Sum2_out6 Sum2_out7 Sum2_out8 Sum2_out9 Sum3_in0 Sum3_in1
+ Sum3_in2 Sum3_in3 Sum3_in4 Sum3_in5 Sum3_in6 Sum3_in7 Sum3_in8 Sum3_in9 Sum3_out0 Sum3_out1
+ Sum3_out2 Sum3_out3 Sum3_out4 Sum3_out5 Sum3_out6 Sum3_out7 Sum3_out8 Sum3_out9 gnd! sel0_reg
+ sel1_reg sel2_reg sel3_reg vdd!
** N=10128 EP=204 FDC=26592
X645 A3_3 A2_3 A1_3 A0_3 B0_reg0 A3_1 gnd! 12 Cin0_3 CLK
+ RST A0_3_8 vdd! A2_1 13 Cin0_2 A0_2_8 A1_1 14 Cin0_1
+ A0_1_8 A0_1 B0_1 60 B0_0 B0_2 B0_3 Cin0_0 A0_0_8 A3_2
+ A2_2 A1_2 A0_2 B0_reg1 9 A3_0 10 A2_0 11 A1_0
+ 52 A0_0 B0_reg2 51 5 4 3 A0_3_9 A0_2_9 A0_1_9
+ A0_0_9 B0_reg3 6 7 8 53 Sel3 Sel2 Sel1 Sel0
+ 30 29 28 27 Sum0_in0 Sum0_in1 Sum0_in2 Sum0_in3 Sum0_in7 Sum0_in4
+ Sum0_in8 Sum0_in5 Sum0_in9 Sum0_in6 Sum0_out0 Sum0_out2 Sum0_out9 Sum0_out1 Sum0_out3 Sum0_out7
+ Sum0_out4 Sum0_out8 Sum0_out5 Sum0_out6 ph2p3_Matrix_vector_Multiplication $T=-650 60 0 0 $X=-390 $Y=0
X646 12 13 14 60 B1_reg0 3 gnd! 24 Cin1_3 CLK
+ RST A1_3_8 vdd! 4 25 Cin1_2 A1_2_8 5 26 Cin1_1
+ A1_1_8 51 B1_1 61 B1_0 B1_2 B1_3 Cin1_0 A1_0_8 9
+ 10 11 52 B1_reg1 21 6 22 7 23 8
+ 55 53 B1_reg2 54 17 16 15 A1_3_9 A1_2_9 A1_1_9
+ A1_0_9 B1_reg3 18 19 20 56 27 28 29 30
+ 46 45 44 43 Sum1_in0 Sum1_in1 Sum1_in2 Sum1_in3 Sum1_in7 Sum1_in4
+ Sum1_in8 Sum1_in5 Sum1_in9 Sum1_in6 Sum1_out0 Sum1_out2 Sum1_out9 Sum1_out1 Sum1_out3 Sum1_out7
+ Sum1_out4 Sum1_out8 Sum1_out5 Sum1_out6 ph2p3_Matrix_vector_Multiplication $T=63440 60 0 0 $X=63700 $Y=0
X647 24 25 26 61 B2_reg0 15 gnd! 40 Cin2_3 CLK
+ RST A2_3_8 vdd! 16 41 Cin2_2 A2_2_8 17 42 Cin2_1
+ A2_1_8 54 B2_1 62 B2_0 B2_2 B2_3 Cin2_0 A2_0_8 21
+ 22 23 55 B2_reg1 37 18 38 19 39 20
+ 58 56 B2_reg2 57 33 32 31 A2_3_9 A2_2_9 A2_1_9
+ A2_0_9 B2_reg3 34 35 36 59 43 44 45 46
+ 50 49 48 47 Sum2_in0 Sum2_in1 Sum2_in2 Sum2_in3 Sum2_in7 Sum2_in4
+ Sum2_in8 Sum2_in5 Sum2_in9 Sum2_in6 Sum2_out0 Sum2_out2 Sum2_out9 Sum2_out1 Sum2_out3 Sum2_out7
+ Sum2_out4 Sum2_out8 Sum2_out5 Sum2_out6 ph2p3_Matrix_vector_Multiplication $T=127530 60 0 0 $X=127790 $Y=0
X648 40 41 42 62 B3_reg0 31 gnd! A3_reg3 Cin3_3 CLK
+ RST A3_3_8 vdd! 32 A2_reg3 Cin3_2 A3_2_8 33 A1_reg3 Cin3_1
+ A3_1_8 57 B3_1 A0_reg3 B3_0 B3_2 B3_3 Cin3_0 A3_0_8 37
+ 38 39 58 B3_reg1 A3_reg2 34 A2_reg2 35 A1_reg2 36
+ A0_reg2 59 B3_reg2 A0_reg1 A1_reg1 A2_reg1 A3_reg1 A3_3_9 A3_2_9 A3_1_9
+ A3_0_9 B3_reg3 A3_reg0 A2_reg0 A1_reg0 A0_reg0 47 48 49 50
+ sel0_reg sel1_reg sel2_reg sel3_reg Sum3_in0 Sum3_in1 Sum3_in2 Sum3_in3 Sum3_in7 Sum3_in4
+ Sum3_in8 Sum3_in5 Sum3_in9 Sum3_in6 Sum3_out0 Sum3_out2 Sum3_out9 Sum3_out1 Sum3_out3 Sum3_out7
+ Sum3_out4 Sum3_out8 Sum3_out5 Sum3_out6 ph2p3_Matrix_vector_Multiplication $T=191620 60 0 0 $X=191880 $Y=0
.ends ph3_sytolic_array
