* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : NAND2_2X                                     *
* Netlisted  : Mon Sep 30 17:00:58 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_3 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 2 3 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=20.4563 scb=0.0180281 scc=0.00115498 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_4 1 2 3 4
** N=4 EP=4 FDC=1
M0 1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_5                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_5 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 3 2 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=24.7379 scb=0.0260985 scc=0.00157851 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_6                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_6 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_2X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_2X 5 1 2 4 3
** N=6 EP=5 FDC=4
X0 1 M1_PO_CDNS_1 $T=520 1760 0 90 $X=400 $Y=1660
X1 2 M1_PO_CDNS_1 $T=1200 1820 0 90 $X=1080 $Y=1720
X2 3 2 4 5 3 pmos1v_CDNS_3 $T=1030 2070 0 0 $X=790 $Y=1870
X3 4 2 6 5 nmos1v_CDNS_4 $T=830 710 0 0 $X=630 $Y=510
X4 4 3 1 5 3 pmos1v_CDNS_5 $T=620 2070 0 0 $X=200 $Y=1870
X5 5 1 6 nmos1v_CDNS_6 $T=620 710 0 0 $X=200 $Y=510
.ends NAND2_2X
