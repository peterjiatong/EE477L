* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 8bit_CSA                                     *
* Netlisted  : Sun Nov  3 07:45:00 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_8                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_8 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_16                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_16 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_18                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_18 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_19                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_19 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR2_1X                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR2_1X 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=10
X0 1 M1_PO_CDNS_8 $T=580 2010 0 90 $X=460 $Y=1910
X1 2 M1_PO_CDNS_8 $T=1490 1580 0 90 $X=1370 $Y=1480
X2 6 M1_PO_CDNS_8 $T=3880 1920 0 90 $X=3760 $Y=1820
X3 7 M1_PO_CDNS_8 $T=4800 1580 0 90 $X=4680 $Y=1480
X4 6 M2_M1_CDNS_16 $T=1040 1920 0 90 $X=910 $Y=1840
X5 7 M2_M1_CDNS_16 $T=1960 1580 0 90 $X=1830 $Y=1500
X6 8 M2_M1_CDNS_16 $T=3270 3070 0 0 $X=3190 $Y=2940
X7 9 M2_M1_CDNS_16 $T=3360 690 0 90 $X=3230 $Y=610
X8 6 M2_M1_CDNS_16 $T=3460 1920 0 90 $X=3330 $Y=1840
X9 8 M2_M1_CDNS_16 $T=3790 3050 0 0 $X=3710 $Y=2920
X10 7 M2_M1_CDNS_16 $T=4520 1580 0 90 $X=4390 $Y=1500
X11 8 M2_M1_CDNS_16 $T=4720 3050 0 0 $X=4640 $Y=2920
X12 9 M2_M1_CDNS_16 $T=5550 690 0 90 $X=5420 $Y=610
X13 8 M2_M1_CDNS_16 $T=5650 3050 0 0 $X=5570 $Y=2920
X14 4 1 6 4 nmos1v_CDNS_18 $T=650 860 0 0 $X=230 $Y=660
X15 4 2 7 4 nmos1v_CDNS_18 $T=1580 860 0 0 $X=1160 $Y=660
X16 4 2 9 4 nmos1v_CDNS_18 $T=3020 860 0 0 $X=2600 $Y=660
X17 10 6 5 4 nmos1v_CDNS_18 $T=3950 860 0 0 $X=3530 $Y=660
X18 10 7 4 4 nmos1v_CDNS_18 $T=4880 860 0 0 $X=4460 $Y=660
X19 9 1 5 4 nmos1v_CDNS_18 $T=5810 860 0 0 $X=5390 $Y=660
X20 3 1 6 4 3 pmos1v_CDNS_19 $T=650 2490 0 0 $X=230 $Y=2290
X21 3 2 7 4 3 pmos1v_CDNS_19 $T=1580 2490 0 0 $X=1160 $Y=2290
X22 3 2 8 4 3 pmos1v_CDNS_19 $T=3020 2500 0 0 $X=2600 $Y=2300
X23 8 6 5 4 3 pmos1v_CDNS_19 $T=3950 2500 0 0 $X=3530 $Y=2300
X24 8 7 5 4 3 pmos1v_CDNS_19 $T=4880 2500 0 0 $X=4460 $Y=2300
X25 8 1 3 4 3 pmos1v_CDNS_19 $T=5810 2500 0 0 $X=5390 $Y=2300
M0 6 1 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=650 $Y=860 $dt=0
M1 7 2 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1580 $Y=860 $dt=0
M2 9 2 4 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=3020 $Y=860 $dt=0
M3 5 6 10 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=3950 $Y=860 $dt=0
M4 4 7 10 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4880 $Y=860 $dt=0
M5 5 1 9 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5810 $Y=860 $dt=0
M6 8 2 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3020 $Y=2500 $dt=1
M7 5 6 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3950 $Y=2500 $dt=1
M8 5 7 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=4880 $Y=2500 $dt=1
M9 3 1 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=5810 $Y=2500 $dt=1
.ends XOR2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_11                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_11 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X 1 2 3 4 5 6
** N=6 EP=6 FDC=4
X0 1 M1_PO_CDNS_8 $T=520 1770 0 90 $X=400 $Y=1670
X1 4 M1_PO_CDNS_8 $T=1200 1830 0 90 $X=1080 $Y=1730
X2 2 3 cellTmpl_CDNS_11 $T=120 150 0 0 $X=0 $Y=10
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=620 $Y=720 $dt=0
M1 5 4 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=830 $Y=720 $dt=0
M2 5 1 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=620 $Y=2080 $dt=1
M3 2 4 5 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=1030 $Y=2080 $dt=1
.ends NAND2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_2X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_2X 1 2 3 4 5 6
** N=6 EP=6 FDC=4
X0 3 M1_PO_CDNS_8 $T=520 1760 0 90 $X=400 $Y=1660
X1 4 M1_PO_CDNS_8 $T=1200 1820 0 90 $X=1080 $Y=1720
X2 1 2 cellTmpl_CDNS_11 $T=120 140 0 0 $X=0 $Y=0
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=620 $Y=710 $dt=0
M1 5 4 6 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=830 $Y=710 $dt=0
M2 5 3 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=15.9511 scb=0.0138709 scc=0.00113792 $X=620 $Y=2070 $dt=1
M3 1 4 5 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=15.9511 scb=0.0138709 scc=0.00113792 $X=1030 $Y=2070 $dt=1
.ends NAND2_2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 1_bit_Full_Adder_ver1                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 1_bit_Full_Adder_ver1 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=23 EP=12 FDC=34
X0 2 M3_M2_CDNS_1 $T=1170 1430 0 0 $X=1090 $Y=1180
X1 3 M3_M2_CDNS_1 $T=8020 1830 0 90 $X=7770 $Y=1750
X2 2 M3_M2_CDNS_1 $T=8650 1560 0 0 $X=8570 $Y=1310
X3 6 M3_M2_CDNS_1 $T=12070 1330 0 0 $X=11990 $Y=1080
X4 3 M3_M2_CDNS_1 $T=12670 2160 0 0 $X=12590 $Y=1910
X5 2 M2_M1_CDNS_2 $T=1170 1430 0 0 $X=1090 $Y=1180
X6 3 M2_M1_CDNS_2 $T=8020 1830 0 90 $X=7770 $Y=1750
X7 2 M2_M1_CDNS_2 $T=8650 1560 0 0 $X=8570 $Y=1310
X8 6 M2_M1_CDNS_2 $T=12070 1330 0 0 $X=11990 $Y=1080
X9 3 M2_M1_CDNS_2 $T=12670 2160 0 0 $X=12590 $Y=1910
X10 1 M4_M3_CDNS_3 $T=270 1810 0 0 $X=190 $Y=1560
X11 8 M4_M3_CDNS_3 $T=6460 1360 0 0 $X=6380 $Y=1110
X12 9 M4_M3_CDNS_3 $T=8070 1290 0 0 $X=7990 $Y=1040
X13 1 M4_M3_CDNS_3 $T=10010 1820 0 90 $X=9760 $Y=1740
X14 9 M4_M3_CDNS_3 $T=12110 1830 0 90 $X=11860 $Y=1750
X15 8 M4_M3_CDNS_3 $T=13590 1430 0 0 $X=13510 $Y=1180
X16 1 M3_M2_CDNS_4 $T=270 1810 0 0 $X=190 $Y=1560
X17 8 M3_M2_CDNS_4 $T=6460 1360 0 0 $X=6380 $Y=1110
X18 9 M3_M2_CDNS_4 $T=8070 1290 0 0 $X=7990 $Y=1040
X19 1 M3_M2_CDNS_4 $T=10010 1820 0 90 $X=9760 $Y=1740
X20 9 M3_M2_CDNS_4 $T=12110 1830 0 90 $X=11860 $Y=1750
X21 8 M3_M2_CDNS_4 $T=13590 1430 0 0 $X=13510 $Y=1180
X22 1 M2_M1_CDNS_5 $T=270 1810 0 0 $X=190 $Y=1560
X23 8 M2_M1_CDNS_5 $T=6460 1360 0 0 $X=6380 $Y=1110
X24 9 M2_M1_CDNS_5 $T=8070 1290 0 0 $X=7990 $Y=1040
X25 1 M2_M1_CDNS_5 $T=10010 1820 0 90 $X=9760 $Y=1740
X26 9 M2_M1_CDNS_5 $T=12110 1830 0 90 $X=11860 $Y=1750
X27 8 M2_M1_CDNS_5 $T=13590 1430 0 0 $X=13510 $Y=1180
X28 2 5 4 1 10 18 NAND2_1X $T=8400 -10 0 0 $X=8400 $Y=0
X29 10 5 4 9 6 19 NAND2_1X $T=10400 -10 0 0 $X=10400 $Y=0
X30 5 4 8 3 9 17 NAND2_2X $T=6400 0 0 0 $X=6400 $Y=0
X31 1 2 5 4 8 11 12 22 15 16 XOR2_1X $T=0 0 0 0 $X=0 $Y=0
X32 3 8 5 4 7 13 14 23 20 21 XOR2_1X $T=12400 0 0 0 $X=12400 $Y=0
M0 13 3 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=13050 $Y=2490 $dt=1
M1 14 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=13980 $Y=2490 $dt=1
.ends 1_bit_Full_Adder_ver1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X 1 2 3 4
** N=4 EP=4 FDC=2
X0 4 M1_PO_CDNS_8 $T=970 1740 0 90 $X=850 $Y=1640
X1 2 3 cellTmpl_CDNS_11 $T=130 140 0 0 $X=10 $Y=0
M0 1 4 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6908 scb=0.0179614 scc=0.00130074 $X=1090 $Y=1110 $dt=0
M1 1 4 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=18.2452 scb=0.0177397 scc=0.00150411 $X=1090 $Y=2120 $dt=1
.ends INV_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND4_1x                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND4_1x 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=15 EP=12 FDC=18
X0 2 3 4 1 8 13 NAND2_1X $T=0 -10 0 0 $X=0 $Y=0
X1 5 3 4 6 9 14 NAND2_1X $T=4000 -10 0 0 $X=4000 $Y=0
X2 10 3 4 11 12 15 NAND2_1X $T=8000 -10 0 0 $X=8000 $Y=0
X3 11 M2_M1_CDNS_16 $T=3610 1720 0 90 $X=3480 $Y=1640
X4 11 M2_M1_CDNS_16 $T=9560 1830 0 90 $X=9430 $Y=1750
X5 11 3 4 8 INV_1X $T=1990 0 0 0 $X=2000 $Y=0
X6 10 3 4 9 INV_1X $T=5990 0 0 0 $X=6000 $Y=0
X7 7 3 4 12 INV_1X $T=9990 0 0 0 $X=10000 $Y=0
.ends AND4_1x

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_1X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_1X 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=12 EP=12 FDC=11
X0 2 M1_PO_CDNS_8 $T=670 1870 0 90 $X=550 $Y=1770
X1 7 M1_PO_CDNS_8 $T=1120 1850 0 90 $X=1000 $Y=1750
X2 4 M1_PO_CDNS_8 $T=3920 1900 0 90 $X=3800 $Y=1800
X3 5 M1_PO_CDNS_8 $T=4860 1910 0 90 $X=4740 $Y=1810
X4 8 M1_PO_CDNS_8 $T=6230 1520 0 90 $X=6110 $Y=1420
X5 9 M2_M1_CDNS_16 $T=2390 1260 0 0 $X=2310 $Y=1130
X6 10 M2_M1_CDNS_16 $T=2390 2860 0 0 $X=2310 $Y=2730
X7 9 M2_M1_CDNS_16 $T=3830 1260 0 0 $X=3750 $Y=1130
X8 10 M2_M1_CDNS_16 $T=4770 2860 0 0 $X=4690 $Y=2730
X9 3 2 7 3 nmos1v_CDNS_18 $T=750 890 0 0 $X=330 $Y=690
X10 3 7 9 3 nmos1v_CDNS_18 $T=2140 890 0 0 $X=1720 $Y=690
X11 3 2 11 3 nmos1v_CDNS_18 $T=3070 890 0 0 $X=2650 $Y=690
X12 9 4 8 3 nmos1v_CDNS_18 $T=4000 890 0 0 $X=3580 $Y=690
X13 11 5 8 3 nmos1v_CDNS_18 $T=4930 890 0 0 $X=4510 $Y=690
X14 3 8 6 3 nmos1v_CDNS_18 $T=6310 890 0 0 $X=5890 $Y=690
X15 1 2 7 3 1 pmos1v_CDNS_19 $T=750 2330 0 0 $X=330 $Y=2130
X16 1 7 10 3 1 pmos1v_CDNS_19 $T=2140 2330 0 0 $X=1720 $Y=2130
X17 1 2 12 3 1 pmos1v_CDNS_19 $T=3070 2330 0 0 $X=2650 $Y=2130
X18 12 4 8 3 1 pmos1v_CDNS_19 $T=4000 2330 0 0 $X=3580 $Y=2130
X19 10 5 8 3 1 pmos1v_CDNS_19 $T=4930 2330 0 0 $X=4510 $Y=2130
X20 1 8 6 3 1 pmos1v_CDNS_19 $T=6310 2330 0 0 $X=5890 $Y=2130
M0 7 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=750 $Y=890 $dt=0
M1 9 7 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=2140 $Y=890 $dt=0
M2 11 2 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=3070 $Y=890 $dt=0
M3 8 4 9 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=4000 $Y=890 $dt=0
M4 8 5 11 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=4930 $Y=890 $dt=0
M5 6 8 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=6310 $Y=890 $dt=0
M6 7 2 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=750 $Y=2330 $dt=1
M7 10 7 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=2140 $Y=2330 $dt=1
M8 12 2 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=3070 $Y=2330 $dt=1
M9 8 4 12 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=4000 $Y=2330 $dt=1
M10 8 5 10 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=4930 $Y=2330 $dt=1
.ends MUX_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CSA                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CSA 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 68
*.DEVICECLIMB
** N=123 EP=28 FDC=219
X0 2 M3_M2_CDNS_1 $T=19990 1430 0 0 $X=19910 $Y=1180
X1 8 M3_M2_CDNS_1 $T=45190 1430 0 0 $X=45110 $Y=1180
X2 11 M3_M2_CDNS_1 $T=70390 1430 0 0 $X=70310 $Y=1180
X3 14 M3_M2_CDNS_1 $T=95590 1430 0 0 $X=95510 $Y=1180
X4 17 M3_M2_CDNS_1 $T=116410 1910 0 0 $X=116330 $Y=1660
X5 3 M3_M2_CDNS_1 $T=117350 2060 0 0 $X=117270 $Y=1810
X6 2 M2_M1_CDNS_2 $T=19990 1430 0 0 $X=19910 $Y=1180
X7 8 M2_M1_CDNS_2 $T=45190 1430 0 0 $X=45110 $Y=1180
X8 11 M2_M1_CDNS_2 $T=70390 1430 0 0 $X=70310 $Y=1180
X9 14 M2_M1_CDNS_2 $T=95590 1430 0 0 $X=95510 $Y=1180
X10 17 M2_M1_CDNS_2 $T=116410 1910 0 0 $X=116330 $Y=1660
X11 3 M2_M1_CDNS_2 $T=117350 2060 0 0 $X=117270 $Y=1810
X12 1 M4_M3_CDNS_3 $T=18950 2010 0 90 $X=18700 $Y=1930
X13 7 M4_M3_CDNS_3 $T=44120 2000 0 90 $X=43870 $Y=1920
X14 10 M4_M3_CDNS_3 $T=69330 2010 0 90 $X=69080 $Y=1930
X15 13 M4_M3_CDNS_3 $T=94500 2000 0 90 $X=94250 $Y=1920
X16 1 M3_M2_CDNS_4 $T=18950 2010 0 90 $X=18700 $Y=1930
X17 18 M3_M2_CDNS_4 $T=24960 1870 0 0 $X=24880 $Y=1620
X18 7 M3_M2_CDNS_4 $T=44120 2000 0 90 $X=43870 $Y=1920
X19 19 M3_M2_CDNS_4 $T=50160 1870 0 0 $X=50080 $Y=1620
X20 10 M3_M2_CDNS_4 $T=69330 2010 0 90 $X=69080 $Y=1930
X21 20 M3_M2_CDNS_4 $T=75360 1870 0 0 $X=75280 $Y=1620
X22 13 M3_M2_CDNS_4 $T=94500 2000 0 90 $X=94250 $Y=1920
X23 20 M3_M2_CDNS_4 $T=102430 1820 0 90 $X=102180 $Y=1740
X24 19 M3_M2_CDNS_4 $T=105050 1610 0 0 $X=104970 $Y=1360
X25 18 M3_M2_CDNS_4 $T=106450 1820 0 90 $X=106200 $Y=1740
X26 1 M2_M1_CDNS_5 $T=18950 2010 0 90 $X=18700 $Y=1930
X27 18 M2_M1_CDNS_5 $T=24960 1870 0 0 $X=24880 $Y=1620
X28 7 M2_M1_CDNS_5 $T=44120 2000 0 90 $X=43870 $Y=1920
X29 19 M2_M1_CDNS_5 $T=50160 1870 0 0 $X=50080 $Y=1620
X30 10 M2_M1_CDNS_5 $T=69330 2010 0 90 $X=69080 $Y=1930
X31 20 M2_M1_CDNS_5 $T=75360 1870 0 0 $X=75280 $Y=1620
X32 13 M2_M1_CDNS_5 $T=94500 2000 0 90 $X=94250 $Y=1920
X33 20 M2_M1_CDNS_5 $T=102430 1820 0 90 $X=102180 $Y=1740
X34 19 M2_M1_CDNS_5 $T=105050 1610 0 0 $X=104970 $Y=1360
X35 18 M2_M1_CDNS_5 $T=106450 1820 0 90 $X=106200 $Y=1740
X36 18 M5_M4_CDNS_6 $T=24960 1870 0 0 $X=24880 $Y=1620
X37 19 M5_M4_CDNS_6 $T=50160 1870 0 0 $X=50080 $Y=1620
X38 20 M5_M4_CDNS_6 $T=75360 1870 0 0 $X=75280 $Y=1620
X39 20 M5_M4_CDNS_6 $T=102430 1820 0 90 $X=102180 $Y=1740
X40 19 M5_M4_CDNS_6 $T=105050 1610 0 0 $X=104970 $Y=1360
X41 18 M5_M4_CDNS_6 $T=106450 1820 0 90 $X=106200 $Y=1740
X42 18 M4_M3_CDNS_7 $T=24960 1870 0 0 $X=24880 $Y=1620
X43 19 M4_M3_CDNS_7 $T=50160 1870 0 0 $X=50080 $Y=1620
X44 20 M4_M3_CDNS_7 $T=75360 1870 0 0 $X=75280 $Y=1620
X45 20 M4_M3_CDNS_7 $T=102430 1820 0 90 $X=102180 $Y=1740
X46 19 M4_M3_CDNS_7 $T=105050 1610 0 0 $X=104970 $Y=1360
X47 18 M4_M3_CDNS_7 $T=106450 1820 0 90 $X=106200 $Y=1740
X48 1 2 4 5 18 33 34 112 76 77 XOR2_1X $T=18800 0 0 0 $X=18800 $Y=0
X49 7 8 4 5 19 42 43 115 85 86 XOR2_1X $T=44000 0 0 0 $X=44000 $Y=0
X50 10 11 4 5 20 51 52 118 94 95 XOR2_1X $T=69200 0 0 0 $X=69200 $Y=0
X51 13 14 4 5 21 60 61 121 103 104 XOR2_1X $T=94400 0 0 0 $X=94400 $Y=0
X52 1 2 3 5 4 22 6 28 30 29
+ 26 27 1_bit_Full_Adder_ver1 $T=0 0 0 0 $X=0 $Y=0
X53 7 8 22 5 4 23 9 37 39 38
+ 35 36 1_bit_Full_Adder_ver1 $T=25200 0 0 0 $X=25200 $Y=0
X54 10 11 23 5 4 24 12 46 48 47
+ 44 45 1_bit_Full_Adder_ver1 $T=50400 0 0 0 $X=50400 $Y=0
X55 13 14 24 5 4 17 15 55 57 56
+ 53 54 1_bit_Full_Adder_ver1 $T=75600 0 0 0 $X=75600 $Y=0
X56 20 21 4 5 19 18 25 62 63 64
+ 65 66 AND4_1x $T=100800 0 0 0 $X=100800 $Y=0
X57 4 25 5 17 3 16 67 68 108 122
+ 109 123 MUX_1X $T=112790 0 0 0 $X=112800 $Y=0
M0 33 1 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=19450 $Y=2490 $dt=1
M1 34 2 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=20380 $Y=2490 $dt=1
M2 35 7 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=25850 $Y=2490 $dt=1
M3 36 8 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=26780 $Y=2490 $dt=1
M4 42 7 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=44650 $Y=2490 $dt=1
M5 43 8 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=45580 $Y=2490 $dt=1
M6 44 10 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=51050 $Y=2490 $dt=1
M7 45 11 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=51980 $Y=2490 $dt=1
M8 51 10 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=69850 $Y=2490 $dt=1
M9 52 11 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=70780 $Y=2490 $dt=1
M10 53 13 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=76250 $Y=2490 $dt=1
M11 54 14 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=77180 $Y=2490 $dt=1
M12 60 13 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=95050 $Y=2490 $dt=1
M13 61 14 4 4 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=95980 $Y=2490 $dt=1
.ends 4bit_CSA

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 8bit_CSA                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 8bit_CSA 2 8 11 14 17 20 23 26 3 9
+ 12 15 18 21 24 27 4 29 7 10
+ 13 16 19 22 25 28 6 5
** N=243 EP=28 FDC=444
X0 1 M3_M2_CDNS_1 $T=119680 1510 0 0 $X=119600 $Y=1260
X1 1 M2_M1_CDNS_2 $T=119680 1510 0 0 $X=119600 $Y=1260
X2 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 1 80 73 72 70
+ 69 42 52 62 79 30 31 81 4bit_CSA $T=0 0 0 0 $X=0 $Y=0
X3 17 18 1 5 6 19 20 21 22 23
+ 24 25 26 27 28 29 132 125 124 122
+ 121 94 104 114 131 82 83 133 4bit_CSA $T=119800 0 0 0 $X=119800 $Y=0
M0 30 2 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=17.6861 scb=0.0184591 scc=0.000433664 $X=650 $Y=2490 $dt=1
M1 31 3 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.886 scb=0.00790338 scc=9.25552e-05 $X=1580 $Y=2490 $dt=1
M2 1 81 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=119100 $Y=2330 $dt=1
M3 82 17 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=120450 $Y=2490 $dt=1
M4 83 18 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=121380 $Y=2490 $dt=1
M5 29 133 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=19.0824 scb=0.0208702 scc=0.000619562 $X=238900 $Y=2330 $dt=1
.ends 8bit_CSA
