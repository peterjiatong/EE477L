* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph1p3_MSDFF                                  *
* Netlisted  : Sat Nov 23 21:33:14 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_8                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_8 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_10                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_10 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_11                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_11 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 1 M1_PO_CDNS_8 $T=700 2040 0 90 $X=580 $Y=1940
X1 3 1 4 3 nmos1v_CDNS_10 $T=780 900 0 0 $X=360 $Y=700
X2 2 4 1 3 2 pmos1v_CDNS_11 $T=780 2430 0 0 $X=360 $Y=2230
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=780 $Y=900 $dt=0
.ends INV_1X_small_layout

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_12                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_12 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_8 $T=640 1830 0 90 $X=520 $Y=1730
X1 6 M1_PO_CDNS_8 $T=1940 640 0 0 $X=1840 $Y=520
X2 3 1 6 3 nmos1v_CDNS_10 $T=710 860 0 0 $X=290 $Y=660
X3 4 6 5 3 nmos1v_CDNS_10 $T=1890 860 0 0 $X=1470 $Y=660
X4 2 3 cellTmpl_CDNS_12 $T=120 140 0 0 $X=0 $Y=0
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=710 $Y=860 $dt=0
M1 5 6 4 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1890 $Y=860 $dt=0
.ends ph1p3_clk_part

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X_small                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X_small 1 2 3 4 5 6
** N=6 EP=6 FDC=4
X0 3 M1_PO_CDNS_8 $T=690 1680 0 90 $X=570 $Y=1580
X1 5 M1_PO_CDNS_8 $T=1930 1650 0 90 $X=1810 $Y=1550
X2 2 3 6 2 nmos1v_CDNS_10 $T=810 1000 0 0 $X=390 $Y=800
X3 6 5 4 2 nmos1v_CDNS_10 $T=2050 1000 0 0 $X=1630 $Y=800
X4 1 4 3 2 1 pmos1v_CDNS_11 $T=810 2440 0 0 $X=390 $Y=2240
X5 1 4 5 2 1 pmos1v_CDNS_11 $T=2050 2450 0 0 $X=1630 $Y=2250
X6 1 2 cellTmpl_CDNS_12 $T=240 210 0 0 $X=120 $Y=70
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=810 $Y=1000 $dt=0
M1 4 5 6 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=2050 $Y=1000 $dt=0
M2 4 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=810 $Y=2440 $dt=1
M3 4 5 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=2050 $Y=2450 $dt=1
.ends NAND2_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_14                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_14 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_MSDFF                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_MSDFF 1 13 4 11 12 10
** N=18 EP=6 FDC=30
X0 1 M2_M1_CDNS_1 $T=430 2010 0 0 $X=350 $Y=1880
X1 2 M2_M1_CDNS_1 $T=1110 -1470 0 0 $X=1030 $Y=-1600
X2 1 M2_M1_CDNS_1 $T=2790 -1820 0 0 $X=2710 $Y=-1950
X3 3 M2_M1_CDNS_1 $T=4150 -1460 0 180 $X=4070 $Y=-1590
X4 4 M2_M1_CDNS_1 $T=5200 -2030 0 0 $X=5120 $Y=-2160
X5 2 M2_M1_CDNS_1 $T=5310 1560 0 90 $X=5180 $Y=1480
X6 3 M2_M1_CDNS_1 $T=5670 -1460 0 90 $X=5540 $Y=-1540
X7 5 M2_M1_CDNS_1 $T=6280 1490 0 0 $X=6200 $Y=1360
X8 6 M2_M1_CDNS_1 $T=7300 1510 0 90 $X=7170 $Y=1430
X9 5 M2_M1_CDNS_1 $T=7850 -2080 0 0 $X=7770 $Y=-2210
X10 6 M2_M1_CDNS_1 $T=9400 1510 0 90 $X=9270 $Y=1430
X11 4 M2_M1_CDNS_1 $T=9770 -2060 0 0 $X=9690 $Y=-2190
X12 7 M3_M2_CDNS_2 $T=1140 2170 0 90 $X=890 $Y=2090
X13 8 M3_M2_CDNS_2 $T=3910 970 0 0 $X=3830 $Y=720
X14 9 M3_M2_CDNS_2 $T=4630 -2070 0 180 $X=4550 $Y=-2320
X15 7 M3_M2_CDNS_2 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X16 7 M3_M2_CDNS_2 $T=8100 2170 0 90 $X=7850 $Y=2090
X17 9 M3_M2_CDNS_2 $T=8890 -1970 0 180 $X=8810 $Y=-2220
X18 8 M3_M2_CDNS_2 $T=9760 1890 0 0 $X=9680 $Y=1640
X19 10 M2_M1_CDNS_3 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X20 10 M2_M1_CDNS_3 $T=5110 3310 0 0 $X=5030 $Y=3060
X21 7 M2_M1_CDNS_3 $T=8100 2170 0 90 $X=7850 $Y=2090
X22 7 M2_M1_CDNS_5 $T=1140 2170 0 90 $X=890 $Y=2090
X23 8 M2_M1_CDNS_5 $T=3910 970 0 0 $X=3830 $Y=720
X24 9 M2_M1_CDNS_5 $T=4630 -2070 0 180 $X=4550 $Y=-2320
X25 7 M2_M1_CDNS_5 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X26 9 M2_M1_CDNS_5 $T=8890 -1970 0 180 $X=8810 $Y=-2220
X27 8 M2_M1_CDNS_5 $T=9760 1890 0 0 $X=9680 $Y=1640
X28 10 M4_M3_CDNS_6 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X29 10 M4_M3_CDNS_6 $T=5110 3310 0 0 $X=5030 $Y=3060
X30 10 M3_M2_CDNS_7 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X31 10 M3_M2_CDNS_7 $T=5110 3310 0 0 $X=5030 $Y=3060
X32 11 10 12 2 INV_1X_small_layout $T=0 40 1 0 $X=0 $Y=-3760
X33 1 10 12 7 INV_1X_small_layout $T=0 0 0 0 $X=0 $Y=0
X34 4 10 12 3 INV_1X_small_layout $T=4800 40 1 0 $X=4800 $Y=-3760
X35 5 10 12 6 INV_1X_small_layout $T=6200 0 0 0 $X=6200 $Y=0
X36 9 10 12 4 INV_1X_small_layout $T=8600 40 1 0 $X=8600 $Y=-3760
X37 1 10 12 13 8 14 ph1p3_clk_part $T=1400 0 0 0 $X=1400 $Y=0
X38 1 10 12 3 9 15 ph1p3_clk_part $T=2400 40 1 0 $X=2400 $Y=-3760
X39 7 10 12 5 9 16 ph1p3_clk_part $T=6200 40 1 0 $X=6200 $Y=-3760
X40 7 10 12 6 8 17 ph1p3_clk_part $T=7600 0 0 0 $X=7600 $Y=0
X41 10 12 8 5 2 18 NAND2_1X_small $T=3680 -70 0 0 $X=3800 $Y=0
X42 10 12 cellTmpl_CDNS_14 $T=1520 -100 1 0 $X=1400 $Y=-3760
M0 2 11 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=780 $Y=-2870 $dt=1
M1 7 1 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=780 $Y=2430 $dt=1
M2 14 1 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=2110 $Y=2460 $dt=1
M3 15 1 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=3110 $Y=-2900 $dt=1
M4 8 1 13 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=3290 $Y=2460 $dt=1
M5 9 1 3 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=4290 $Y=-2660 $dt=1
M6 3 4 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=5580 $Y=-2870 $dt=1
M7 16 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=6910 $Y=-2900 $dt=1
M8 6 5 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=6980 $Y=2430 $dt=1
M9 9 7 5 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=8090 $Y=-2660 $dt=1
M10 17 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=8310 $Y=2460 $dt=1
M11 4 9 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=9380 $Y=-2870 $dt=1
M12 8 7 6 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=9490 $Y=2460 $dt=1
.ends ph1p3_MSDFF
