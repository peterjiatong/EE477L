* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : INV_2X                                       *
* Netlisted  : Mon Sep 30 15:08:49 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_3 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 1 3 2 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.0576 scb=0.0170651 scc=0.000872115 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_4 1 2 3
** N=3 EP=3 FDC=1
M0 1 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=17.8161 scb=0.0190899 scc=0.00152594 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_2X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_2X 4 3 1 2
** N=4 EP=4 FDC=2
X0 1 2 3 4 2 pmos1v_CDNS_3 $T=1030 2110 0 0 $X=610 $Y=1910
X1 1 4 3 nmos1v_CDNS_4 $T=1030 1130 0 0 $X=610 $Y=930
.ends INV_2X
