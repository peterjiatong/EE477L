* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph2p3_Matrix_vector_Multiplication           *
* Netlisted  : Tue Dec  3 19:35:00 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_8                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_8 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_9                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_9 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_10                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_10 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_11                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_11 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_12                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_12 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_13                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_13 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_14                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_14 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_15                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_15 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_16                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_16 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_17                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_17 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_18                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_18 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_new                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_new 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 3 M1_PO_CDNS_16 $T=1020 1750 0 90 $X=900 $Y=1650
X1 1 2 cellTmpl_CDNS_18 $T=50 150 0 0 $X=-70 $Y=10
M0 4 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.3086 scb=0.00950139 scc=0.000267597 $X=1140 $Y=930 $dt=0
.ends INV_1X_new

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_19                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_19 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_20                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_20 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_20

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_21                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_21 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_21

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X_small                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_16 $T=690 1680 0 90 $X=570 $Y=1580
X1 4 M1_PO_CDNS_16 $T=1930 1650 0 90 $X=1810 $Y=1550
X2 3 1 6 3 nmos1v_CDNS_19 $T=810 1000 0 0 $X=390 $Y=800
X3 6 4 5 3 nmos1v_CDNS_19 $T=2050 1000 0 0 $X=1630 $Y=800
X4 2 1 5 3 2 pmos1v_CDNS_20 $T=810 2440 0 0 $X=390 $Y=2240
X5 2 4 5 3 2 pmos1v_CDNS_20 $T=2050 2450 0 0 $X=1630 $Y=2250
X6 2 3 cellTmpl_CDNS_21 $T=240 210 0 0 $X=120 $Y=70
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=810 $Y=1000 $dt=0
M1 5 4 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=2050 $Y=1000 $dt=0
.ends NAND2_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6
*.DEVICECLIMB
** N=7 EP=6 FDC=3
X0 2 3 6 5 INV_1X_new $T=2480 -10 0 0 $X=2410 $Y=0
X1 1 2 3 4 6 7 NAND2_1X_small $T=-110 -70 0 0 $X=10 $Y=0
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_22                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_22 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_23                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_23 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_23

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_24                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_24 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_24

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_25                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_25 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_25

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_26                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_26 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_26

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_27                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_27 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_27

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_28                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_28 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_28

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_29                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_29 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_29

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR_small                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR_small 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=9
X0 1 M2_M1_CDNS_11 $T=350 1340 0 90 $X=220 $Y=1260
X1 6 M2_M1_CDNS_11 $T=5510 3180 0 90 $X=5380 $Y=3100
X2 6 M2_M1_CDNS_11 $T=6740 3180 0 90 $X=6610 $Y=3100
X3 1 M1_PO_CDNS_16 $T=580 1660 0 90 $X=460 $Y=1560
X4 4 M1_PO_CDNS_16 $T=1990 1480 0 90 $X=1870 $Y=1380
X5 4 M1_PO_CDNS_22 $T=5990 1680 0 90 $X=5790 $Y=1580
X6 1 M1_PO_CDNS_22 $T=7100 1350 0 90 $X=6900 $Y=1250
X7 7 M1_PO_CDNS_23 $T=3070 1660 0 90 $X=2870 $Y=1560
X8 8 M1_PO_CDNS_23 $T=4410 1540 0 90 $X=4210 $Y=1440
X9 8 M3_M2_CDNS_24 $T=1210 1540 0 90 $X=1010 $Y=1440
X10 8 M3_M2_CDNS_24 $T=4410 1540 0 90 $X=4210 $Y=1440
X11 8 M2_M1_CDNS_25 $T=1210 1540 0 90 $X=1010 $Y=1440
X12 4 M2_M1_CDNS_25 $T=1820 1880 0 90 $X=1620 $Y=1780
X13 8 M2_M1_CDNS_25 $T=4410 1540 0 90 $X=4210 $Y=1440
X14 4 M2_M1_CDNS_26 $T=5990 1680 0 90 $X=5790 $Y=1580
X15 1 M2_M1_CDNS_26 $T=7100 1350 0 90 $X=6900 $Y=1250
X16 2 3 cellTmpl_CDNS_27 $T=120 140 0 0 $X=0 $Y=0
X17 2 1 8 3 2 pmos1v_CDNS_28 $T=700 2180 0 0 $X=280 $Y=1980
X18 2 4 7 3 2 pmos1v_CDNS_28 $T=2110 2170 0 0 $X=1690 $Y=1970
X19 2 7 6 3 2 pmos1v_CDNS_28 $T=3270 2160 0 0 $X=2850 $Y=1960
X20 2 8 6 3 2 pmos1v_CDNS_28 $T=4610 2160 0 0 $X=4190 $Y=1960
X21 6 4 5 3 2 pmos1v_CDNS_28 $T=6140 2120 0 0 $X=5720 $Y=1920
X22 6 1 5 3 2 pmos1v_CDNS_28 $T=7250 2160 0 0 $X=6830 $Y=1960
X23 3 1 8 3 nmos1v_CDNS_29 $T=700 590 0 0 $X=280 $Y=390
X24 3 4 7 3 nmos1v_CDNS_29 $T=2110 580 0 0 $X=1690 $Y=380
X25 3 7 9 3 nmos1v_CDNS_29 $T=3270 580 0 0 $X=2850 $Y=380
X26 9 8 5 3 nmos1v_CDNS_29 $T=4610 580 0 0 $X=4190 $Y=380
X27 3 4 10 3 nmos1v_CDNS_29 $T=6140 600 0 0 $X=5720 $Y=400
X28 10 1 5 3 nmos1v_CDNS_29 $T=7250 650 0 0 $X=6830 $Y=450
M0 8 1 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.45462 scb=0.00478425 scc=6.8709e-05 $X=700 $Y=590 $dt=0
M1 7 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=2110 $Y=580 $dt=0
M2 9 7 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=3270 $Y=580 $dt=0
M3 5 8 9 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=4610 $Y=580 $dt=0
M4 10 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 $X=6140 $Y=600 $dt=0
M5 5 1 10 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=7250 $Y=650 $dt=0
M6 7 4 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.1869 scb=0.0086398 scc=0.00051649 $X=2110 $Y=2170 $dt=1
M7 6 7 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3270 $Y=2160 $dt=1
M8 6 8 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4610 $Y=2160 $dt=1
.ends XOR_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 8 9 13
*.DEVICECLIMB
** N=13 EP=9 FDC=12
X0 4 M3_M2_CDNS_1 $T=6750 2480 0 0 $X=6670 $Y=2230
X1 4 M3_M2_CDNS_1 $T=9120 2880 0 0 $X=9040 $Y=2630
X2 4 M2_M1_CDNS_10 $T=6750 2480 0 0 $X=6670 $Y=2230
X3 4 M2_M1_CDNS_10 $T=9120 2880 0 0 $X=9040 $Y=2630
X4 4 M1_PO_CDNS_13 $T=6750 2480 0 0 $X=6650 $Y=2230
X5 4 M1_PO_CDNS_13 $T=9120 2880 0 0 $X=9020 $Y=2630
X6 1 3 2 4 6 9 AND $T=7790 0 0 0 $X=7800 $Y=0
X7 1 3 2 4 5 13 7 8 10 11 XOR_small $T=0 0 0 0 $X=0 $Y=0
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_33                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_33 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_33

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_1X_small                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=-310 120 0 0 $X=-430 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1000 $Y=830 $dt=0
M1 4 5 6 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1210 $Y=830 $dt=0
.ends NAND_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_2X_small1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_2X_small1 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=130 160 0 0 $X=10 $Y=20
M0 6 4 2 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=7.66878 scb=0.00580736 scc=7.77234e-05 $X=940 $Y=890 $dt=0
M1 3 5 6 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=11.676 scb=0.0124835 scc=0.000479408 $X=940 $Y=1100 $dt=0
.ends NAND_2X_small1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_39                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_39 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_39

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR1 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=6
X0 6 M2_M1_CDNS_11 $T=1210 1480 0 90 $X=1080 $Y=1400
X1 7 M2_M1_CDNS_11 $T=2250 1860 0 90 $X=2120 $Y=1780
X2 6 M2_M1_CDNS_11 $T=2950 1480 0 90 $X=2820 $Y=1400
X3 8 M2_M1_CDNS_11 $T=3370 650 0 0 $X=3290 $Y=520
X4 9 M2_M1_CDNS_11 $T=3370 3080 0 0 $X=3290 $Y=2950
X5 9 M2_M1_CDNS_11 $T=3930 3080 0 0 $X=3850 $Y=2950
X6 7 M2_M1_CDNS_11 $T=4680 1860 0 90 $X=4550 $Y=1780
X7 9 M2_M1_CDNS_11 $T=4890 3070 0 0 $X=4810 $Y=2940
X8 8 M2_M1_CDNS_11 $T=5840 640 0 0 $X=5760 $Y=510
X9 9 M2_M1_CDNS_11 $T=6260 3080 0 0 $X=6180 $Y=2950
X10 6 M1_PO_CDNS_16 $T=4020 1500 0 90 $X=3900 $Y=1400
X11 7 M1_PO_CDNS_16 $T=5020 1730 0 90 $X=4900 $Y=1630
X12 2 3 6 2 nmos1v_CDNS_19 $T=830 840 0 0 $X=410 $Y=640
X13 2 4 7 2 nmos1v_CDNS_19 $T=1790 840 0 0 $X=1370 $Y=640
X14 1 3 6 2 1 pmos1v_CDNS_20 $T=830 2320 0 0 $X=410 $Y=2120
X15 1 4 7 2 1 pmos1v_CDNS_20 $T=1790 2320 0 0 $X=1370 $Y=2120
X16 1 4 9 2 1 pmos1v_CDNS_28 $T=3120 2080 0 0 $X=2700 $Y=1880
X17 9 6 5 2 1 pmos1v_CDNS_28 $T=4090 2140 0 0 $X=3670 $Y=1940
X18 9 7 5 2 1 pmos1v_CDNS_28 $T=5050 2140 0 0 $X=4630 $Y=1940
X19 1 3 9 2 1 pmos1v_CDNS_28 $T=6010 2140 0 0 $X=5590 $Y=1940
X20 2 4 8 2 nmos1v_CDNS_29 $T=3120 780 0 0 $X=2700 $Y=580
X21 10 6 5 2 nmos1v_CDNS_29 $T=4090 760 0 0 $X=3670 $Y=560
X22 10 7 2 2 nmos1v_CDNS_29 $T=5050 770 0 0 $X=4630 $Y=570
X23 8 3 5 2 nmos1v_CDNS_29 $T=6010 770 0 0 $X=5590 $Y=570
X24 1 2 cellTmpl_CDNS_39 $T=180 120 0 0 $X=60 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=830 $Y=840 $dt=0
M1 7 4 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1790 $Y=840 $dt=0
M2 8 4 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=3120 $Y=780 $dt=0
M3 5 6 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4126 scb=0.0095497 scc=0.000351079 $X=4090 $Y=760 $dt=0
M4 2 7 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=5050 $Y=770 $dt=0
M5 5 3 8 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=6010 $Y=770 $dt=0
.ends XOR1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder1_small                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder1_small 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 22 23
*.DEVICECLIMB
** N=23 EP=16 FDC=18
X0 1 M3_M2_CDNS_1 $T=590 2080 0 90 $X=340 $Y=2000
X1 3 M3_M2_CDNS_1 $T=2300 3150 0 90 $X=2050 $Y=3070
X2 1 M3_M2_CDNS_1 $T=17380 1890 0 0 $X=17300 $Y=1640
X3 3 M3_M2_CDNS_1 $T=19040 3010 0 0 $X=18960 $Y=2760
X4 1 M2_M1_CDNS_10 $T=590 2080 0 90 $X=340 $Y=2000
X5 3 M2_M1_CDNS_10 $T=2300 3150 0 90 $X=2050 $Y=3070
X6 1 M2_M1_CDNS_10 $T=17380 1890 0 0 $X=17300 $Y=1640
X7 3 M2_M1_CDNS_10 $T=19040 3010 0 0 $X=18960 $Y=2760
X8 8 M2_M1_CDNS_11 $T=6580 1900 0 0 $X=6500 $Y=1770
X9 9 M2_M1_CDNS_11 $T=15190 1730 0 90 $X=15060 $Y=1650
X10 1 M1_PO_CDNS_13 $T=590 2080 0 90 $X=340 $Y=1980
X11 3 M1_PO_CDNS_13 $T=2300 3150 0 90 $X=2050 $Y=3050
X12 1 M1_PO_CDNS_13 $T=17380 1890 0 0 $X=17280 $Y=1640
X13 3 M1_PO_CDNS_13 $T=19040 3010 0 0 $X=18940 $Y=2760
X14 8 M3_M2_CDNS_14 $T=6970 950 0 0 $X=6890 $Y=820
X15 8 M3_M2_CDNS_14 $T=14100 570 0 90 $X=13970 $Y=490
X16 8 M1_PO_CDNS_15 $T=8510 1970 0 0 $X=8410 $Y=1720
X17 8 M1_PO_CDNS_15 $T=16110 1570 0 0 $X=16010 $Y=1320
X18 9 M1_PO_CDNS_15 $T=20260 1840 0 0 $X=20160 $Y=1590
X19 1 M1_PO_CDNS_16 $T=690 1610 0 0 $X=590 $Y=1490
X20 3 M1_PO_CDNS_16 $T=1650 1990 0 0 $X=1550 $Y=1870
X21 5 M1_PO_CDNS_16 $T=7590 1960 0 0 $X=7490 $Y=1840
X22 10 M1_PO_CDNS_16 $T=19320 1680 0 0 $X=19220 $Y=1560
X23 8 M2_M1_CDNS_17 $T=8510 1970 0 0 $X=8430 $Y=1720
X24 8 M2_M1_CDNS_17 $T=16110 1570 0 0 $X=16030 $Y=1320
X25 9 M2_M1_CDNS_17 $T=20260 1840 0 0 $X=20180 $Y=1590
X26 2 4 1 10 3 20 NAND_1X_small $T=16970 30 0 0 $X=16540 $Y=10
X27 2 4 9 7 10 21 NAND_1X_small $T=19810 30 0 0 $X=19380 $Y=10
X28 2 4 9 5 8 19 NAND_2X_small1 $T=13690 -10 0 0 $X=13700 $Y=10
X29 2 4 1 3 8 11 12 15 22 16 XOR1 $T=-40 30 0 0 $X=20 $Y=10
X30 2 4 5 8 6 13 14 17 23 18 XOR1 $T=6800 30 0 0 $X=6860 $Y=10
.ends full_adder1_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: multiplier                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt multiplier 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
** N=238 EP=50 FDC=456
X0 2 M3_M2_CDNS_1 $T=160 15480 0 0 $X=80 $Y=15230
X1 2 M3_M2_CDNS_1 $T=160 21130 0 0 $X=80 $Y=20880
X2 2 M3_M2_CDNS_1 $T=170 9270 0 0 $X=90 $Y=9020
X3 2 M3_M2_CDNS_1 $T=170 13790 0 0 $X=90 $Y=13540
X4 19 M3_M2_CDNS_1 $T=500 8210 0 0 $X=420 $Y=7960
X5 1 M3_M2_CDNS_1 $T=1350 15570 0 0 $X=1270 $Y=15320
X6 1 M3_M2_CDNS_1 $T=1360 13320 0 0 $X=1280 $Y=13070
X7 20 M3_M2_CDNS_1 $T=4380 23070 0 90 $X=4130 $Y=22990
X8 21 M3_M2_CDNS_1 $T=4340 15320 0 0 $X=4260 $Y=15070
X9 22 M3_M2_CDNS_1 $T=5400 21130 0 0 $X=5320 $Y=20880
X10 7 M3_M2_CDNS_1 $T=5740 15570 0 0 $X=5660 $Y=15320
X11 7 M3_M2_CDNS_1 $T=5750 13320 0 0 $X=5670 $Y=13070
X12 19 M3_M2_CDNS_1 $T=6590 5910 0 0 $X=6510 $Y=5660
X13 23 M3_M2_CDNS_1 $T=7520 22860 0 0 $X=7440 $Y=22610
X14 23 M3_M2_CDNS_1 $T=7960 21030 0 0 $X=7880 $Y=20780
X15 24 M3_M2_CDNS_1 $T=8730 15340 0 0 $X=8650 $Y=15090
X16 8 M3_M2_CDNS_1 $T=8980 17010 0 0 $X=8900 $Y=16760
X17 8 M3_M2_CDNS_1 $T=10140 15570 0 0 $X=10060 $Y=15320
X18 8 M3_M2_CDNS_1 $T=10150 13320 0 0 $X=10070 $Y=13070
X19 25 M3_M2_CDNS_1 $T=12100 19160 0 0 $X=12020 $Y=18910
X20 20 M3_M2_CDNS_1 $T=12260 20780 0 0 $X=12180 $Y=20530
X21 26 M3_M2_CDNS_1 $T=13150 15340 0 0 $X=13070 $Y=15090
X22 27 M3_M2_CDNS_1 $T=14690 20780 0 0 $X=14610 $Y=20530
X23 28 M3_M2_CDNS_1 $T=15670 8330 0 0 $X=15590 $Y=8080
X24 29 M3_M2_CDNS_1 $T=16600 750 0 0 $X=16520 $Y=500
X25 27 M3_M2_CDNS_1 $T=17570 22850 0 0 $X=17490 $Y=22600
X26 30 M3_M2_CDNS_1 $T=22230 22840 0 0 $X=22150 $Y=22590
X27 30 M3_M2_CDNS_1 $T=28820 20830 0 0 $X=28740 $Y=20580
X28 31 M3_M2_CDNS_1 $T=35370 22940 0 0 $X=35290 $Y=22690
X29 2 M2_M1_CDNS_2 $T=160 15480 0 0 $X=80 $Y=15230
X30 2 M2_M1_CDNS_2 $T=160 21130 0 0 $X=80 $Y=20880
X31 2 M2_M1_CDNS_2 $T=170 9270 0 0 $X=90 $Y=9020
X32 2 M2_M1_CDNS_2 $T=170 13790 0 0 $X=90 $Y=13540
X33 19 M2_M1_CDNS_2 $T=500 8210 0 0 $X=420 $Y=7960
X34 20 M2_M1_CDNS_2 $T=4380 23070 0 90 $X=4130 $Y=22990
X35 21 M2_M1_CDNS_2 $T=4340 15320 0 0 $X=4260 $Y=15070
X36 22 M2_M1_CDNS_2 $T=5400 21130 0 0 $X=5320 $Y=20880
X37 24 M2_M1_CDNS_2 $T=8730 15340 0 0 $X=8650 $Y=15090
X38 25 M2_M1_CDNS_2 $T=12100 19160 0 0 $X=12020 $Y=18910
X39 26 M2_M1_CDNS_2 $T=13150 15340 0 0 $X=13070 $Y=15090
X40 27 M2_M1_CDNS_2 $T=17570 22850 0 0 $X=17490 $Y=22600
X41 30 M2_M1_CDNS_2 $T=22230 22840 0 0 $X=22150 $Y=22590
X42 30 M2_M1_CDNS_2 $T=28820 20830 0 0 $X=28740 $Y=20580
X43 31 M2_M1_CDNS_2 $T=35370 22940 0 0 $X=35290 $Y=22690
X44 32 M2_M1_CDNS_2 $T=46340 18970 0 0 $X=46260 $Y=18720
X45 30 M5_M4_CDNS_3 $T=28820 19250 0 0 $X=28740 $Y=19120
X46 33 M5_M4_CDNS_3 $T=35550 19590 0 0 $X=35470 $Y=19460
X47 1 M3_M2_CDNS_4 $T=1390 19500 0 0 $X=1310 $Y=19250
X48 21 M3_M2_CDNS_4 $T=3370 8280 0 0 $X=3290 $Y=8030
X49 34 M3_M2_CDNS_4 $T=5400 9800 0 0 $X=5320 $Y=9550
X50 7 M3_M2_CDNS_4 $T=7950 19550 0 0 $X=7870 $Y=19300
X51 25 M3_M2_CDNS_4 $T=12950 9830 0 0 $X=12870 $Y=9580
X52 35 M3_M2_CDNS_4 $T=14070 2580 0 90 $X=13820 $Y=2500
X53 36 M3_M2_CDNS_4 $T=15700 9710 0 0 $X=15620 $Y=9460
X54 11 M3_M2_CDNS_4 $T=25590 19380 0 0 $X=25510 $Y=19130
X55 37 M3_M2_CDNS_4 $T=25970 20660 0 0 $X=25890 $Y=20410
X56 38 M3_M2_CDNS_4 $T=28540 8430 0 0 $X=28460 $Y=8180
X57 38 M3_M2_CDNS_4 $T=28700 9810 0 0 $X=28620 $Y=9560
X58 32 M3_M2_CDNS_4 $T=38260 18710 0 0 $X=38180 $Y=18460
X59 39 M3_M2_CDNS_4 $T=42090 2930 0 90 $X=41840 $Y=2850
X60 30 M4_M3_CDNS_5 $T=28820 19250 0 0 $X=28740 $Y=19000
X61 30 M4_M3_CDNS_5 $T=34220 19150 0 0 $X=34140 $Y=18900
X62 1 M4_M3_CDNS_6 $T=1390 19500 0 0 $X=1310 $Y=19250
X63 21 M4_M3_CDNS_6 $T=3370 8280 0 0 $X=3290 $Y=8030
X64 7 M4_M3_CDNS_6 $T=4510 16920 0 0 $X=4430 $Y=16670
X65 34 M4_M3_CDNS_6 $T=5400 9800 0 0 $X=5320 $Y=9550
X66 7 M4_M3_CDNS_6 $T=7950 19550 0 0 $X=7870 $Y=19300
X67 40 M4_M3_CDNS_6 $T=8750 8160 0 0 $X=8670 $Y=7910
X68 41 M4_M3_CDNS_6 $T=10750 19470 0 0 $X=10670 $Y=19220
X69 42 M4_M3_CDNS_6 $T=11680 11800 0 0 $X=11600 $Y=11550
X70 25 M4_M3_CDNS_6 $T=12950 9830 0 0 $X=12870 $Y=9580
X71 11 M4_M3_CDNS_6 $T=13290 16990 0 0 $X=13210 $Y=16740
X72 35 M4_M3_CDNS_6 $T=14070 2580 0 90 $X=13820 $Y=2500
X73 36 M4_M3_CDNS_6 $T=15700 9710 0 0 $X=15620 $Y=9460
X74 42 M4_M3_CDNS_6 $T=22150 6400 0 0 $X=22070 $Y=6150
X75 36 M4_M3_CDNS_6 $T=24490 750 0 0 $X=24410 $Y=500
X76 11 M4_M3_CDNS_6 $T=25590 19380 0 0 $X=25510 $Y=19130
X77 37 M4_M3_CDNS_6 $T=25970 20660 0 0 $X=25890 $Y=20410
X78 43 M4_M3_CDNS_6 $T=26370 19410 0 0 $X=26290 $Y=19160
X79 33 M4_M3_CDNS_6 $T=26600 23000 0 0 $X=26520 $Y=22750
X80 38 M4_M3_CDNS_6 $T=28540 8430 0 0 $X=28460 $Y=8180
X81 38 M4_M3_CDNS_6 $T=28700 9810 0 0 $X=28620 $Y=9560
X82 44 M4_M3_CDNS_6 $T=29280 19170 0 0 $X=29200 $Y=18920
X83 39 M4_M3_CDNS_6 $T=35970 2380 0 0 $X=35890 $Y=2130
X84 32 M4_M3_CDNS_6 $T=38260 18710 0 0 $X=38180 $Y=18460
X85 44 M4_M3_CDNS_6 $T=39640 17490 0 0 $X=39560 $Y=17240
X86 39 M4_M3_CDNS_6 $T=42090 2930 0 90 $X=41840 $Y=2850
X87 28 M4_M3_CDNS_6 $T=43850 8260 0 0 $X=43770 $Y=8010
X88 29 M4_M3_CDNS_6 $T=43880 660 0 0 $X=43800 $Y=410
X89 32 M4_M3_CDNS_6 $T=46340 18970 0 0 $X=46260 $Y=18720
X90 30 M5_M4_CDNS_7 $T=34220 19150 0 0 $X=34140 $Y=18900
X91 33 M5_M4_CDNS_7 $T=34850 16990 0 0 $X=34770 $Y=16740
X92 1 M4_M3_CDNS_8 $T=1390 21140 0 0 $X=1310 $Y=21010
X93 21 M4_M3_CDNS_8 $T=3650 6110 0 0 $X=3570 $Y=5980
X94 34 M4_M3_CDNS_8 $T=6680 2460 0 0 $X=6600 $Y=2330
X95 37 M4_M3_CDNS_8 $T=13170 22790 0 0 $X=13090 $Y=22660
X96 25 M4_M3_CDNS_8 $T=13680 4950 0 0 $X=13600 $Y=4820
X97 11 M4_M3_CDNS_8 $T=14530 13310 0 0 $X=14450 $Y=13180
X98 11 M4_M3_CDNS_8 $T=14530 15600 0 0 $X=14450 $Y=15470
X99 35 M4_M3_CDNS_8 $T=21870 1570 0 0 $X=21790 $Y=1440
X100 40 M4_M3_CDNS_8 $T=23120 3950 0 0 $X=23040 $Y=3820
X101 43 M4_M3_CDNS_8 $T=28320 12210 0 0 $X=28240 $Y=12080
X102 29 M4_M3_CDNS_8 $T=28540 230 0 90 $X=28410 $Y=150
X103 28 M4_M3_CDNS_8 $T=28550 7610 0 90 $X=28420 $Y=7530
X104 41 M4_M3_CDNS_8 $T=33860 19960 0 90 $X=33730 $Y=19880
X105 1 M3_M2_CDNS_9 $T=1390 21140 0 0 $X=1310 $Y=20890
X106 7 M3_M2_CDNS_9 $T=4510 16920 0 0 $X=4430 $Y=16670
X107 40 M3_M2_CDNS_9 $T=8750 8160 0 0 $X=8670 $Y=7910
X108 41 M3_M2_CDNS_9 $T=10750 19470 0 0 $X=10670 $Y=19220
X109 42 M3_M2_CDNS_9 $T=11680 11800 0 0 $X=11600 $Y=11550
X110 37 M3_M2_CDNS_9 $T=13170 22790 0 0 $X=13090 $Y=22540
X111 11 M3_M2_CDNS_9 $T=13290 16990 0 0 $X=13210 $Y=16740
X112 11 M3_M2_CDNS_9 $T=14530 13310 0 0 $X=14450 $Y=13060
X113 11 M3_M2_CDNS_9 $T=14530 15600 0 0 $X=14450 $Y=15350
X114 42 M3_M2_CDNS_9 $T=22150 6400 0 0 $X=22070 $Y=6150
X115 36 M3_M2_CDNS_9 $T=24490 750 0 0 $X=24410 $Y=500
X116 43 M3_M2_CDNS_9 $T=26370 19410 0 0 $X=26290 $Y=19160
X117 33 M3_M2_CDNS_9 $T=26600 23000 0 0 $X=26520 $Y=22750
X118 30 M3_M2_CDNS_9 $T=28820 19250 0 0 $X=28740 $Y=19000
X119 44 M3_M2_CDNS_9 $T=29280 19170 0 0 $X=29200 $Y=18920
X120 41 M3_M2_CDNS_9 $T=33860 19960 0 90 $X=33610 $Y=19880
X121 30 M3_M2_CDNS_9 $T=34220 19150 0 0 $X=34140 $Y=18900
X122 39 M3_M2_CDNS_9 $T=35970 2380 0 0 $X=35890 $Y=2130
X123 44 M3_M2_CDNS_9 $T=39640 17490 0 0 $X=39560 $Y=17240
X124 28 M3_M2_CDNS_9 $T=43850 8260 0 0 $X=43770 $Y=8010
X125 29 M3_M2_CDNS_9 $T=43880 660 0 0 $X=43800 $Y=410
X126 32 M3_M2_CDNS_9 $T=46340 18970 0 0 $X=46260 $Y=18720
X127 1 M2_M1_CDNS_10 $T=1350 15570 0 0 $X=1270 $Y=15320
X128 1 M2_M1_CDNS_10 $T=1360 13320 0 0 $X=1280 $Y=13070
X129 1 M2_M1_CDNS_10 $T=1390 21140 0 0 $X=1310 $Y=20890
X130 7 M2_M1_CDNS_10 $T=4510 16920 0 0 $X=4430 $Y=16670
X131 7 M2_M1_CDNS_10 $T=5740 15570 0 0 $X=5660 $Y=15320
X132 7 M2_M1_CDNS_10 $T=5750 13320 0 0 $X=5670 $Y=13070
X133 19 M2_M1_CDNS_10 $T=6590 5910 0 0 $X=6510 $Y=5660
X134 23 M2_M1_CDNS_10 $T=7520 22860 0 0 $X=7440 $Y=22610
X135 23 M2_M1_CDNS_10 $T=7960 21030 0 0 $X=7880 $Y=20780
X136 40 M2_M1_CDNS_10 $T=8750 8160 0 0 $X=8670 $Y=7910
X137 8 M2_M1_CDNS_10 $T=8980 17010 0 0 $X=8900 $Y=16760
X138 8 M2_M1_CDNS_10 $T=10140 15570 0 0 $X=10060 $Y=15320
X139 8 M2_M1_CDNS_10 $T=10150 13320 0 0 $X=10070 $Y=13070
X140 8 M2_M1_CDNS_10 $T=10370 18740 0 0 $X=10290 $Y=18490
X141 41 M2_M1_CDNS_10 $T=10750 19470 0 0 $X=10670 $Y=19220
X142 42 M2_M1_CDNS_10 $T=11680 11800 0 0 $X=11600 $Y=11550
X143 20 M2_M1_CDNS_10 $T=12260 20780 0 0 $X=12180 $Y=20530
X144 37 M2_M1_CDNS_10 $T=13170 22790 0 0 $X=13090 $Y=22540
X145 11 M2_M1_CDNS_10 $T=13290 16990 0 0 $X=13210 $Y=16740
X146 11 M2_M1_CDNS_10 $T=14530 13310 0 0 $X=14450 $Y=13060
X147 11 M2_M1_CDNS_10 $T=14530 15600 0 0 $X=14450 $Y=15350
X148 27 M2_M1_CDNS_10 $T=14690 20780 0 0 $X=14610 $Y=20530
X149 28 M2_M1_CDNS_10 $T=15670 8330 0 0 $X=15590 $Y=8080
X150 29 M2_M1_CDNS_10 $T=16600 750 0 0 $X=16520 $Y=500
X151 42 M2_M1_CDNS_10 $T=22150 6400 0 0 $X=22070 $Y=6150
X152 36 M2_M1_CDNS_10 $T=24490 750 0 0 $X=24410 $Y=500
X153 43 M2_M1_CDNS_10 $T=26370 19410 0 0 $X=26290 $Y=19160
X154 33 M2_M1_CDNS_10 $T=26600 23000 0 0 $X=26520 $Y=22750
X155 30 M2_M1_CDNS_10 $T=28820 19250 0 0 $X=28740 $Y=19000
X156 44 M2_M1_CDNS_10 $T=29280 19170 0 0 $X=29200 $Y=18920
X157 41 M2_M1_CDNS_10 $T=33860 19960 0 90 $X=33610 $Y=19880
X158 30 M2_M1_CDNS_10 $T=34220 19150 0 0 $X=34140 $Y=18900
X159 31 M2_M1_CDNS_10 $T=35760 21100 0 0 $X=35680 $Y=20850
X160 39 M2_M1_CDNS_10 $T=35970 2380 0 0 $X=35890 $Y=2130
X161 44 M2_M1_CDNS_10 $T=39640 17490 0 0 $X=39560 $Y=17240
X162 28 M2_M1_CDNS_10 $T=43850 8260 0 0 $X=43770 $Y=8010
X163 29 M2_M1_CDNS_10 $T=43880 660 0 0 $X=43800 $Y=410
X164 2 M2_M1_CDNS_11 $T=170 4730 0 0 $X=90 $Y=4600
X165 2 M2_M1_CDNS_11 $T=180 890 0 0 $X=100 $Y=760
X166 34 M2_M1_CDNS_11 $T=4340 11800 0 0 $X=4260 $Y=11670
X167 36 M2_M1_CDNS_11 $T=8880 12210 0 0 $X=8800 $Y=12080
X168 35 M2_M1_CDNS_11 $T=13420 4530 0 0 $X=13340 $Y=4400
X169 45 M2_M1_CDNS_11 $T=17560 15460 0 0 $X=17480 $Y=15330
X170 46 M2_M1_CDNS_11 $T=21930 4780 0 0 $X=21850 $Y=4650
X171 38 M2_M1_CDNS_11 $T=29730 11900 0 0 $X=29650 $Y=11770
X172 47 M2_M1_CDNS_11 $T=31310 15530 0 0 $X=31230 $Y=15400
X173 48 M2_M1_CDNS_11 $T=35410 9580 0 0 $X=35330 $Y=9450
X174 49 M2_M1_CDNS_11 $T=41980 11840 0 0 $X=41900 $Y=11710
X175 39 M2_M1_CDNS_11 $T=43890 4790 0 0 $X=43810 $Y=4660
X176 33 M4_M3_CDNS_12 $T=34850 16990 0 0 $X=34770 $Y=16740
X177 1 M1_PO_CDNS_13 $T=1350 15570 0 0 $X=1250 $Y=15320
X178 1 M1_PO_CDNS_13 $T=1360 13320 0 0 $X=1260 $Y=13070
X179 7 M1_PO_CDNS_13 $T=4510 16920 0 0 $X=4410 $Y=16670
X180 7 M1_PO_CDNS_13 $T=5740 15570 0 0 $X=5640 $Y=15320
X181 7 M1_PO_CDNS_13 $T=5750 13320 0 0 $X=5650 $Y=13070
X182 19 M1_PO_CDNS_13 $T=6590 5910 0 0 $X=6490 $Y=5660
X183 23 M1_PO_CDNS_13 $T=7520 22860 0 0 $X=7420 $Y=22610
X184 23 M1_PO_CDNS_13 $T=7960 21030 0 0 $X=7860 $Y=20780
X185 8 M1_PO_CDNS_13 $T=8980 17010 0 0 $X=8880 $Y=16760
X186 8 M1_PO_CDNS_13 $T=10140 15570 0 0 $X=10040 $Y=15320
X187 8 M1_PO_CDNS_13 $T=10150 13320 0 0 $X=10050 $Y=13070
X188 8 M1_PO_CDNS_13 $T=10370 18740 0 0 $X=10270 $Y=18490
X189 41 M1_PO_CDNS_13 $T=10750 19470 0 0 $X=10650 $Y=19220
X190 20 M1_PO_CDNS_13 $T=12260 20780 0 0 $X=12160 $Y=20530
X191 11 M1_PO_CDNS_13 $T=13290 16990 0 0 $X=13190 $Y=16740
X192 11 M1_PO_CDNS_13 $T=14530 13310 0 0 $X=14430 $Y=13060
X193 11 M1_PO_CDNS_13 $T=14530 15600 0 0 $X=14430 $Y=15350
X194 27 M1_PO_CDNS_13 $T=14690 20780 0 0 $X=14590 $Y=20530
X195 28 M1_PO_CDNS_13 $T=15670 8330 0 0 $X=15570 $Y=8080
X196 29 M1_PO_CDNS_13 $T=16600 750 0 0 $X=16500 $Y=500
X197 42 M1_PO_CDNS_13 $T=22150 6400 0 0 $X=22050 $Y=6150
X198 36 M1_PO_CDNS_13 $T=24490 750 0 0 $X=24390 $Y=500
X199 44 M1_PO_CDNS_13 $T=29280 19170 0 0 $X=29180 $Y=18920
X200 30 M1_PO_CDNS_13 $T=34220 19150 0 0 $X=34120 $Y=18900
X201 31 M1_PO_CDNS_13 $T=35760 21100 0 0 $X=35660 $Y=20850
X202 39 M1_PO_CDNS_13 $T=35970 2380 0 0 $X=35870 $Y=2130
X203 21 M3_M2_CDNS_14 $T=4340 13390 0 0 $X=4260 $Y=13260
X204 22 M3_M2_CDNS_14 $T=7370 12440 0 0 $X=7290 $Y=12310
X205 22 M3_M2_CDNS_14 $T=8600 9080 0 0 $X=8520 $Y=8950
X206 8 M3_M2_CDNS_14 $T=10370 18740 0 0 $X=10290 $Y=18610
X207 25 M3_M2_CDNS_14 $T=13190 12020 0 0 $X=13110 $Y=11890
X208 46 M3_M2_CDNS_14 $T=19690 2880 0 90 $X=19560 $Y=2800
X209 37 M3_M2_CDNS_14 $T=26840 17540 0 90 $X=26710 $Y=17460
X210 31 M3_M2_CDNS_14 $T=35760 21100 0 0 $X=35680 $Y=20970
X211 1 M1_PO_CDNS_15 $T=1390 17230 0 0 $X=1290 $Y=16980
X212 1 M1_PO_CDNS_15 $T=1390 24660 0 0 $X=1290 $Y=24410
X213 3 M1_PO_CDNS_15 $T=2770 22320 0 90 $X=2520 $Y=22220
X214 5 M1_PO_CDNS_15 $T=2650 13610 0 0 $X=2550 $Y=13360
X215 4 M1_PO_CDNS_15 $T=2750 17050 0 0 $X=2650 $Y=16800
X216 1 M1_PO_CDNS_15 $T=4410 23850 0 0 $X=4310 $Y=23600
X217 4 M1_PO_CDNS_15 $T=5790 16970 0 0 $X=5690 $Y=16720
X218 9 M1_PO_CDNS_15 $T=7290 23970 0 90 $X=7040 $Y=23870
X219 5 M1_PO_CDNS_15 $T=7180 13450 0 0 $X=7080 $Y=13200
X220 3 M1_PO_CDNS_15 $T=8720 22330 0 90 $X=8470 $Y=22230
X221 3 M1_PO_CDNS_15 $T=9910 24890 0 90 $X=9660 $Y=24790
X222 4 M1_PO_CDNS_15 $T=10210 17010 0 0 $X=10110 $Y=16760
X223 7 M1_PO_CDNS_15 $T=11550 22710 0 0 $X=11450 $Y=22460
X224 5 M1_PO_CDNS_15 $T=11730 13390 0 0 $X=11630 $Y=13140
X225 9 M1_PO_CDNS_15 $T=13230 23970 0 90 $X=12980 $Y=23870
X226 4 M1_PO_CDNS_15 $T=14630 17040 0 0 $X=14530 $Y=16790
X227 7 M1_PO_CDNS_15 $T=15790 22330 0 90 $X=15540 $Y=22230
X228 5 M1_PO_CDNS_15 $T=15980 13520 0 0 $X=15880 $Y=13270
X229 3 M1_PO_CDNS_15 $T=17780 24480 0 0 $X=17680 $Y=24230
X230 8 M1_PO_CDNS_15 $T=20560 22320 0 90 $X=20310 $Y=22220
X231 9 M1_PO_CDNS_15 $T=22240 23950 0 0 $X=22140 $Y=23700
X232 8 M1_PO_CDNS_15 $T=24880 22320 0 90 $X=24630 $Y=22220
X233 3 M1_PO_CDNS_15 $T=26710 24400 0 0 $X=26610 $Y=24150
X234 38 M1_PO_CDNS_15 $T=28540 6330 0 0 $X=28440 $Y=6080
X235 11 M1_PO_CDNS_15 $T=29350 22530 0 0 $X=29250 $Y=22280
X236 45 M1_PO_CDNS_15 $T=29800 13490 0 0 $X=29700 $Y=13240
X237 9 M1_PO_CDNS_15 $T=31140 23850 0 0 $X=31040 $Y=23600
X238 47 M1_PO_CDNS_15 $T=31170 13680 0 0 $X=31070 $Y=13430
X239 32 M1_PO_CDNS_15 $T=31860 16950 0 0 $X=31760 $Y=16700
X240 11 M1_PO_CDNS_15 $T=33650 22300 0 90 $X=33400 $Y=22200
X241 49 M1_PO_CDNS_15 $T=35890 9730 0 0 $X=35790 $Y=9480
X242 1 M2_M1_CDNS_17 $T=1390 17230 0 0 $X=1310 $Y=16980
X243 1 M2_M1_CDNS_17 $T=1390 24660 0 0 $X=1310 $Y=24410
X244 3 M2_M1_CDNS_17 $T=2770 22320 0 90 $X=2520 $Y=22240
X245 5 M2_M1_CDNS_17 $T=2650 13610 0 0 $X=2570 $Y=13360
X246 4 M2_M1_CDNS_17 $T=2750 17050 0 0 $X=2670 $Y=16800
X247 1 M2_M1_CDNS_17 $T=4410 23850 0 0 $X=4330 $Y=23600
X248 4 M2_M1_CDNS_17 $T=5790 16970 0 0 $X=5710 $Y=16720
X249 9 M2_M1_CDNS_17 $T=7290 23970 0 90 $X=7040 $Y=23890
X250 5 M2_M1_CDNS_17 $T=7180 13450 0 0 $X=7100 $Y=13200
X251 3 M2_M1_CDNS_17 $T=8720 22330 0 90 $X=8470 $Y=22250
X252 3 M2_M1_CDNS_17 $T=9910 24890 0 90 $X=9660 $Y=24810
X253 4 M2_M1_CDNS_17 $T=10210 17010 0 0 $X=10130 $Y=16760
X254 7 M2_M1_CDNS_17 $T=11550 22710 0 0 $X=11470 $Y=22460
X255 5 M2_M1_CDNS_17 $T=11730 13390 0 0 $X=11650 $Y=13140
X256 9 M2_M1_CDNS_17 $T=13230 23970 0 90 $X=12980 $Y=23890
X257 4 M2_M1_CDNS_17 $T=14630 17040 0 0 $X=14550 $Y=16790
X258 7 M2_M1_CDNS_17 $T=15790 22330 0 90 $X=15540 $Y=22250
X259 5 M2_M1_CDNS_17 $T=15980 13520 0 0 $X=15900 $Y=13270
X260 3 M2_M1_CDNS_17 $T=17780 24480 0 0 $X=17700 $Y=24230
X261 8 M2_M1_CDNS_17 $T=20560 22320 0 90 $X=20310 $Y=22240
X262 9 M2_M1_CDNS_17 $T=22240 23950 0 0 $X=22160 $Y=23700
X263 8 M2_M1_CDNS_17 $T=24880 22320 0 90 $X=24630 $Y=22240
X264 3 M2_M1_CDNS_17 $T=26710 24400 0 0 $X=26630 $Y=24150
X265 38 M2_M1_CDNS_17 $T=28540 6330 0 0 $X=28460 $Y=6080
X266 11 M2_M1_CDNS_17 $T=29350 22530 0 0 $X=29270 $Y=22280
X267 45 M2_M1_CDNS_17 $T=29800 13490 0 0 $X=29720 $Y=13240
X268 9 M2_M1_CDNS_17 $T=31140 23850 0 0 $X=31060 $Y=23600
X269 47 M2_M1_CDNS_17 $T=31170 13680 0 0 $X=31090 $Y=13430
X270 32 M2_M1_CDNS_17 $T=31860 16950 0 0 $X=31780 $Y=16700
X271 11 M2_M1_CDNS_17 $T=33650 22300 0 90 $X=33400 $Y=22220
X272 49 M2_M1_CDNS_17 $T=35890 9730 0 0 $X=35810 $Y=9480
X273 1 6 2 5 34 77 AND $T=40 14460 1 0 $X=50 $Y=10660
X274 1 6 2 4 21 76 AND $T=40 14420 0 0 $X=50 $Y=14420
X275 1 6 2 3 20 75 AND $T=40 21740 0 0 $X=50 $Y=21740
X276 7 6 2 5 36 80 AND $T=4440 14460 1 0 $X=4450 $Y=10660
X277 7 6 2 4 24 79 AND $T=4440 14420 0 0 $X=4450 $Y=14420
X278 1 6 2 9 23 78 AND $T=4440 21740 0 0 $X=4450 $Y=21740
X279 8 6 2 5 42 83 AND $T=8840 14460 1 0 $X=8850 $Y=10660
X280 8 6 2 4 26 82 AND $T=8840 14420 0 0 $X=8850 $Y=14420
X281 3 6 2 7 37 81 AND $T=8840 21740 0 0 $X=8850 $Y=21740
X282 11 6 2 5 50 93 AND $T=13240 14460 1 0 $X=13250 $Y=10660
X283 11 6 2 4 45 92 AND $T=13240 14420 0 0 $X=13250 $Y=14420
X284 9 6 2 7 27 91 AND $T=13240 21740 0 0 $X=13250 $Y=21740
X285 3 6 2 8 30 104 AND $T=17880 21740 0 0 $X=17890 $Y=21740
X286 9 6 2 8 33 126 AND $T=22280 21740 0 0 $X=22290 $Y=21740
X287 3 6 2 11 14 127 AND $T=26680 21740 0 0 $X=26690 $Y=21740
X288 9 6 2 11 31 131 AND $T=31080 21740 0 0 $X=31090 $Y=21740
X289 23 2 6 41 22 25 73 74 225 half_adder $T=50 21780 1 0 $X=50 $Y=17980
X290 50 2 6 48 13 38 102 103 228 half_adder $T=17640 14460 1 0 $X=17640 $Y=10660
X291 45 2 6 47 17 49 129 130 237 half_adder $T=29830 14460 1 0 $X=29830 $Y=10660
X292 30 2 6 31 18 32 133 134 238 half_adder $T=34210 21780 1 0 $X=34210 $Y=17980
X293 22 6 24 2 28 40 19 67 70 71
+ 65 66 68 69 223 224 full_adder1_small $T=22270 7090 1 180 $X=20 $Y=7100
X294 34 6 46 2 29 10 12 60 63 64
+ 58 59 61 62 221 222 full_adder1_small $T=30 -230 0 0 $X=50 $Y=-220
X295 21 6 25 2 19 35 46 53 56 57
+ 51 52 54 55 219 220 full_adder1_small $T=30 7150 1 0 $X=50 $Y=3340
X296 20 6 27 2 44 43 41 86 89 90
+ 84 85 87 88 226 227 full_adder1_small $T=12230 21790 1 0 $X=12250 $Y=17980
X297 33 6 37 2 32 47 44 96 99 100
+ 94 95 97 98 229 230 full_adder1_small $T=17850 14410 0 0 $X=17870 $Y=14420
X298 36 6 35 2 39 15 29 121 124 125
+ 119 120 122 123 235 236 full_adder1_small $T=21990 -230 0 0 $X=22010 $Y=-220
X299 42 6 40 2 38 16 39 114 117 118
+ 112 113 115 116 233 234 full_adder1_small $T=21990 7150 1 0 $X=22010 $Y=3340
X300 26 6 43 2 49 48 28 107 110 111
+ 105 106 108 109 231 232 full_adder1_small $T=21990 7090 0 0 $X=22010 $Y=7100
M0 77 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=11610 $dt=1
M1 76 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=16790 $dt=1
M2 75 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=24110 $dt=1
M3 73 23 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=16.2188 scb=0.0173423 scc=0.000698846 $X=750 $Y=18640 $dt=1
M4 58 34 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=2120 $dt=1
M5 51 21 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=4320 $dt=1
M6 19 71 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=1070 $Y=9450 $dt=1
M7 6 70 19 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=1480 $Y=9450 $dt=1
M8 59 46 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=2120 $dt=1
M9 52 25 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=4320 $dt=1
M10 77 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=11600 $dt=1
M11 76 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=16800 $dt=1
M12 75 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=24120 $dt=1
M13 221 46 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=1880 $dt=1
M14 219 25 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=4080 $dt=1
M15 34 77 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=11580 $dt=1
M16 21 76 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=16820 $dt=1
M17 20 75 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=24140 $dt=1
M18 71 24 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=3910 $Y=9450 $dt=1
M19 60 58 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=1940 $dt=1
M20 53 51 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=4020 $dt=1
M21 6 22 71 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=4320 $Y=9450 $dt=1
M22 60 59 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=1940 $dt=1
M23 53 52 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=4020 $dt=1
M24 80 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=11610 $dt=1
M25 79 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=16790 $dt=1
M26 78 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=24110 $dt=1
M27 221 34 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=1940 $dt=1
M28 219 21 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=4020 $dt=1
M29 22 41 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=6190 $Y=18700 $dt=1
M30 80 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=11600 $dt=1
M31 79 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=16800 $dt=1
M32 78 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=24120 $dt=1
M33 70 67 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=6890 $Y=9230 $dt=1
M34 6 28 70 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=7300 $Y=9230 $dt=1
M35 22 23 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=7300 $Y=18660 $dt=1
M36 61 29 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=2120 $dt=1
M37 54 19 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=4320 $dt=1
M38 36 80 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=11580 $dt=1
M39 24 79 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=16820 $dt=1
M40 23 78 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=24140 $dt=1
M41 74 23 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=8540 $Y=18930 $dt=1
M42 62 60 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=2120 $dt=1
M43 55 53 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=4320 $dt=1
M44 6 28 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=9370 $Y=9260 $dt=1
M45 83 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=11610 $dt=1
M46 82 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=16790 $dt=1
M47 81 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=24110 $dt=1
M48 74 41 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=9780 $Y=18920 $dt=1
M49 222 60 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=1880 $dt=1
M50 220 53 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=4080 $dt=1
M51 224 69 40 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10330 $Y=9260 $dt=1
M52 83 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=11600 $dt=1
M53 82 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=16800 $dt=1
M54 81 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=24120 $dt=1
M55 10 61 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=1940 $dt=1
M56 35 54 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=4020 $dt=1
M57 224 68 40 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11290 $Y=9260 $dt=1
M58 25 74 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=11460 $Y=18900 $dt=1
M59 10 62 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=1940 $dt=1
M60 35 55 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=4020 $dt=1
M61 6 67 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=12260 $Y=9200 $dt=1
M62 42 83 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=11580 $dt=1
M63 26 82 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=16820 $dt=1
M64 37 81 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=24140 $dt=1
M65 222 29 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=1940 $dt=1
M66 220 19 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=4020 $dt=1
M67 84 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13020 $Y=18960 $dt=1
M68 6 67 69 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13590 $Y=9440 $dt=1
M69 93 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=11610 $dt=1
M70 92 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=16790 $dt=1
M71 91 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=24110 $dt=1
M72 85 27 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13980 $Y=18960 $dt=1
M73 6 28 68 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=14550 $Y=9440 $dt=1
M74 63 29 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=1910 $dt=1
M75 56 19 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=4050 $dt=1
M76 93 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=11600 $dt=1
M77 92 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=16800 $dt=1
M78 91 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=24120 $dt=1
M79 226 27 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=15310 $Y=18720 $dt=1
M80 6 60 63 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=1910 $dt=1
M81 6 53 56 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=4050 $dt=1
M82 6 22 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16210 $Y=9260 $dt=1
M83 86 84 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16280 $Y=18660 $dt=1
M84 50 93 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=11580 $dt=1
M85 45 92 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=16820 $dt=1
M86 27 91 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=24140 $dt=1
M87 223 66 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17170 $Y=9260 $dt=1
M88 86 85 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17240 $Y=18660 $dt=1
M89 64 34 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=2130 $dt=1
M90 57 21 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=4310 $dt=1
M91 223 65 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18130 $Y=9260 $dt=1
M92 226 20 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18200 $Y=18660 $dt=1
M93 6 46 64 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=2130 $dt=1
M94 6 25 57 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=4310 $dt=1
M95 102 50 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=18340 $Y=11320 $dt=1
M96 104 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=18580 $Y=24110 $dt=1
M97 94 33 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=18640 $Y=16760 $dt=1
M98 6 24 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=19100 $Y=9200 $dt=1
M99 95 37 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19600 $Y=16760 $dt=1
M100 104 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=19820 $Y=24120 $dt=1
M101 87 44 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19860 $Y=18960 $dt=1
M102 6 24 66 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20430 $Y=9440 $dt=1
M103 12 63 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=2130 $dt=1
M104 46 56 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=4310 $dt=1
M105 88 86 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20820 $Y=18960 $dt=1
M106 229 37 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=20930 $Y=16520 $dt=1
M107 6 64 12 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=2130 $dt=1
M108 6 57 46 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=4310 $dt=1
M109 6 22 65 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=21390 $Y=9440 $dt=1
M110 30 104 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=21500 $Y=24140 $dt=1
M111 96 94 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=21900 $Y=16580 $dt=1
M112 227 86 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=22150 $Y=18720 $dt=1
M113 119 36 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=2120 $dt=1
M114 112 42 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=4320 $dt=1
M115 105 26 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=9440 $dt=1
M116 96 95 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=22860 $Y=16580 $dt=1
M117 126 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=22980 $Y=24110 $dt=1
M118 43 87 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23120 $Y=18660 $dt=1
M119 120 35 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=2120 $dt=1
M120 113 40 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=4320 $dt=1
M121 106 43 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=9440 $dt=1
M122 13 48 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=23780 $Y=11380 $dt=1
M123 229 33 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23820 $Y=16580 $dt=1
M124 43 88 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24080 $Y=18660 $dt=1
M125 126 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=24220 $Y=24120 $dt=1
M126 13 50 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24890 $Y=11340 $dt=1
M127 227 44 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=25040 $Y=18660 $dt=1
M128 235 35 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=1880 $dt=1
M129 233 40 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=4080 $dt=1
M130 231 43 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=9200 $dt=1
M131 97 32 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=25480 $Y=16760 $dt=1
M132 33 126 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=25900 $Y=24140 $dt=1
M133 121 119 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=1940 $dt=1
M134 114 112 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=4020 $dt=1
M135 107 105 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=9260 $dt=1
M136 103 50 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26130 $Y=11610 $dt=1
M137 98 96 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=26440 $Y=16760 $dt=1
M138 121 120 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=1940 $dt=1
M139 114 113 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=4020 $dt=1
M140 107 106 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=9260 $dt=1
M141 89 44 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27110 $Y=18690 $dt=1
M142 103 48 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27370 $Y=11600 $dt=1
M143 127 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=27380 $Y=24110 $dt=1
M144 6 86 89 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27520 $Y=18690 $dt=1
M145 230 96 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=27770 $Y=16520 $dt=1
M146 235 36 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=1940 $dt=1
M147 233 42 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=4020 $dt=1
M148 231 26 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=9260 $dt=1
M149 127 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=28620 $Y=24120 $dt=1
M150 47 97 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28740 $Y=16580 $dt=1
M151 38 103 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=29050 $Y=11580 $dt=1
M152 122 39 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=2120 $dt=1
M153 115 38 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=4320 $dt=1
M154 108 49 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=9440 $dt=1
M155 47 98 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=29700 $Y=16580 $dt=1
M156 90 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30090 $Y=18950 $dt=1
M157 14 127 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=30300 $Y=24140 $dt=1
M158 6 27 90 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30500 $Y=18950 $dt=1
M159 129 45 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=30530 $Y=11320 $dt=1
M160 123 121 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=2120 $dt=1
M161 116 114 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=4320 $dt=1
M162 109 107 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=9440 $dt=1
M163 230 32 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=30660 $Y=16580 $dt=1
M164 131 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=31780 $Y=24110 $dt=1
M165 236 121 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=1880 $dt=1
M166 234 114 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=4080 $dt=1
M167 232 107 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=9200 $dt=1
M168 99 32 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=32730 $Y=16550 $dt=1
M169 15 122 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=1940 $dt=1
M170 16 115 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=4020 $dt=1
M171 48 108 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=9260 $dt=1
M172 41 89 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=32930 $Y=18950 $dt=1
M173 131 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=33020 $Y=24120 $dt=1
M174 6 96 99 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=33140 $Y=16550 $dt=1
M175 6 90 41 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=33340 $Y=18950 $dt=1
M176 15 123 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=1940 $dt=1
M177 16 116 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=4020 $dt=1
M178 48 109 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=9260 $dt=1
M179 31 131 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=34700 $Y=24140 $dt=1
M180 236 39 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=1940 $dt=1
M181 234 38 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=4020 $dt=1
M182 232 49 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=9260 $dt=1
M183 133 30 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=34910 $Y=18640 $dt=1
M184 100 33 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=35710 $Y=16770 $dt=1
M185 17 47 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=35970 $Y=11380 $dt=1
M186 6 37 100 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=36120 $Y=16770 $dt=1
M187 124 39 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=1910 $dt=1
M188 117 38 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=4050 $dt=1
M189 110 49 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=9230 $dt=1
M190 17 45 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=37080 $Y=11340 $dt=1
M191 6 121 124 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=1910 $dt=1
M192 6 114 117 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=4050 $dt=1
M193 6 107 110 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=9230 $dt=1
M194 130 45 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=38320 $Y=11610 $dt=1
M195 44 99 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=38550 $Y=16770 $dt=1
M196 6 100 44 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=38960 $Y=16770 $dt=1
M197 130 47 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=39560 $Y=11600 $dt=1
M198 125 36 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=2130 $dt=1
M199 118 42 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=4310 $dt=1
M200 111 26 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=9450 $dt=1
M201 6 35 125 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=2130 $dt=1
M202 6 40 118 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=4310 $dt=1
M203 6 43 111 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=9450 $dt=1
M204 18 31 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.2705 scb=0.0126902 scc=0.000796523 $X=40350 $Y=18700 $dt=1
M205 49 130 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=41240 $Y=11580 $dt=1
M206 18 30 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=41460 $Y=18660 $dt=1
M207 29 124 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=2130 $dt=1
M208 39 117 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=4310 $dt=1
M209 28 110 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=42690 $Y=9450 $dt=1
M210 134 30 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42700 $Y=18930 $dt=1
M211 6 125 29 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=2130 $dt=1
M212 6 118 39 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=4310 $dt=1
M213 6 111 28 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=43100 $Y=9450 $dt=1
M214 134 31 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43940 $Y=18920 $dt=1
M215 32 134 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=45620 $Y=18900 $dt=1
.ends multiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_31                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_31 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_31

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_32                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_32 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_32

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_43                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_43 1 2 3 5 6 8
*.DEVICECLIMB
** N=14 EP=6 FDC=2
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=810 $Y=710 $dt=0
M1 8 6 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=4640 $Y=580 $dt=0
.ends cellTmpl_CDNS_43

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_44                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_44 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_44

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_45                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_45 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_45

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=12
X0 7 M3_M2_CDNS_1 $T=250 -3000 0 0 $X=170 $Y=-3250
X1 7 M3_M2_CDNS_1 $T=960 -2040 0 0 $X=880 $Y=-2290
X2 7 M3_M2_CDNS_1 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X3 7 M2_M1_CDNS_2 $T=960 -2040 0 0 $X=880 $Y=-2290
X4 7 M2_M1_CDNS_10 $T=250 -3000 0 0 $X=170 $Y=-3250
X5 7 M2_M1_CDNS_10 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X6 7 M1_PO_CDNS_13 $T=250 -3000 0 0 $X=150 $Y=-3250
X7 7 M1_PO_CDNS_13 $T=2620 -2730 0 0 $X=2520 $Y=-2980
X8 1 M1_PO_CDNS_15 $T=1300 -3500 0 0 $X=1200 $Y=-3750
X9 1 M1_PO_CDNS_15 $T=2660 -4240 0 0 $X=2560 $Y=-4490
X10 1 M1_PO_CDNS_16 $T=680 -3550 0 0 $X=580 $Y=-3670
X11 2 M1_PO_CDNS_16 $T=1300 -2090 0 0 $X=1200 $Y=-2210
X12 5 M1_PO_CDNS_16 $T=4040 -3180 0 0 $X=3940 $Y=-3300
X13 8 M1_PO_CDNS_16 $T=4300 -3670 0 90 $X=4180 $Y=-3770
X14 1 M2_M1_CDNS_17 $T=1300 -3500 0 0 $X=1220 $Y=-3750
X15 1 M2_M1_CDNS_17 $T=2660 -4240 0 0 $X=2580 $Y=-4490
X16 4 7 9 4 nmos1v_CDNS_31 $T=1990 -4420 0 0 $X=1790 $Y=-4620
X17 8 5 10 4 nmos1v_CDNS_31 $T=3370 -4430 0 0 $X=3170 $Y=-4630
X18 8 2 9 4 nmos1v_CDNS_32 $T=1780 -4420 0 0 $X=1360 $Y=-4620
X19 4 1 10 4 nmos1v_CDNS_32 $T=3160 -4430 0 0 $X=2740 $Y=-4630
X20 3 4 1 7 8 6 cellTmpl_CDNS_43 $T=-60 -5080 0 0 $X=-180 $Y=-5220
X21 3 1 11 4 3 pmos1v_CDNS_44 $T=1990 -3120 0 0 $X=1790 $Y=-3320
X22 8 5 12 4 3 pmos1v_CDNS_44 $T=3370 -3190 0 0 $X=3170 $Y=-3390
X23 8 2 11 4 3 pmos1v_CDNS_45 $T=1780 -3120 0 0 $X=1360 $Y=-3320
X24 3 7 12 4 3 pmos1v_CDNS_45 $T=3160 -3190 0 0 $X=2740 $Y=-3390
M0 9 2 8 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1780 $Y=-4420 $dt=0
M1 4 7 9 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1990 $Y=-4420 $dt=0
M2 10 1 4 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3160 $Y=-4430 $dt=0
M3 8 5 10 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3370 $Y=-4430 $dt=0
M4 7 1 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=750 $Y=-2850 $dt=1
M5 11 2 8 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1780 $Y=-3120 $dt=1
M6 3 1 11 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1990 $Y=-3120 $dt=1
M7 12 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3160 $Y=-3190 $dt=1
M8 8 5 12 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3370 $Y=-3190 $dt=1
M9 6 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.2373 scb=0.0194294 scc=0.00149528 $X=4580 $Y=-3180 $dt=1
.ends MUX_2to1___2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FA_4bit                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FA_4bit 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19
** N=83 EP=19 FDC=144
X0 17 M3_M2_CDNS_1 $T=18840 8310 0 0 $X=18760 $Y=8060
X1 18 M3_M2_CDNS_4 $T=19730 4760 0 0 $X=19650 $Y=4510
X2 18 M4_M3_CDNS_6 $T=14030 6120 0 0 $X=13950 $Y=5870
X3 19 M4_M3_CDNS_6 $T=16960 11880 0 0 $X=16880 $Y=11630
X4 18 M4_M3_CDNS_6 $T=19730 4760 0 0 $X=19650 $Y=4510
X5 19 M4_M3_CDNS_6 $T=22610 11350 0 0 $X=22530 $Y=11100
X6 18 M3_M2_CDNS_9 $T=14030 6120 0 0 $X=13950 $Y=5870
X7 19 M3_M2_CDNS_9 $T=16960 11880 0 0 $X=16880 $Y=11630
X8 19 M3_M2_CDNS_9 $T=22610 11350 0 0 $X=22530 $Y=11100
X9 18 M2_M1_CDNS_10 $T=14030 6120 0 0 $X=13950 $Y=5870
X10 19 M2_M1_CDNS_10 $T=16960 11880 0 0 $X=16880 $Y=11630
X11 17 M2_M1_CDNS_10 $T=18840 8310 0 0 $X=18760 $Y=8060
X12 19 M2_M1_CDNS_10 $T=22610 11350 0 0 $X=22530 $Y=11100
X13 5 M2_M1_CDNS_11 $T=-80 3540 0 0 $X=-160 $Y=3410
X14 5 M2_M1_CDNS_11 $T=-80 10890 0 0 $X=-160 $Y=10760
X15 18 M2_M1_CDNS_11 $T=21770 2020 0 0 $X=21690 $Y=1890
X16 17 M2_M1_CDNS_11 $T=21770 5100 0 0 $X=21690 $Y=4970
X17 18 M1_PO_CDNS_13 $T=14030 6120 0 0 $X=13930 $Y=5870
X18 19 M1_PO_CDNS_13 $T=16960 11880 0 0 $X=16860 $Y=11630
X19 17 M1_PO_CDNS_13 $T=18840 8310 0 0 $X=18740 $Y=8060
X20 17 M3_M2_CDNS_14 $T=21980 9220 0 0 $X=21900 $Y=9090
X21 6 5 1 7 11 12 18 43 46 47
+ 41 42 44 45 82 83 full_adder1_small $T=-90 -130 0 0 $X=-70 $Y=-120
X22 8 5 2 7 18 13 17 36 39 40
+ 34 35 37 38 80 81 full_adder1_small $T=-90 7250 1 0 $X=-70 $Y=3440
X23 9 5 3 7 17 14 19 29 32 33
+ 27 28 30 31 78 79 full_adder1_small $T=-90 7190 0 0 $X=-70 $Y=7200
X24 10 5 4 7 19 15 16 22 25 26
+ 20 21 23 24 76 77 full_adder1_small $T=-90 14570 1 0 $X=-70 $Y=10760
M0 41 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=2220 $dt=1
M1 34 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=4420 $dt=1
M2 27 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=9540 $dt=1
M3 20 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=11740 $dt=1
M4 42 1 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=2220 $dt=1
M5 35 2 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=4420 $dt=1
M6 28 3 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=9540 $dt=1
M7 21 4 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=11740 $dt=1
M8 82 1 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=1980 $dt=1
M9 80 2 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=4180 $dt=1
M10 78 3 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=9300 $dt=1
M11 76 4 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=11500 $dt=1
M12 43 41 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=2040 $dt=1
M13 36 34 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=4120 $dt=1
M14 29 27 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=9360 $dt=1
M15 22 20 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=11440 $dt=1
M16 43 42 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=2040 $dt=1
M17 36 35 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=4120 $dt=1
M18 29 28 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=9360 $dt=1
M19 22 21 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=11440 $dt=1
M20 82 6 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=2040 $dt=1
M21 80 8 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=4120 $dt=1
M22 78 9 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=9360 $dt=1
M23 76 10 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=11440 $dt=1
M24 44 11 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=2220 $dt=1
M25 37 18 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=4420 $dt=1
M26 30 17 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=9540 $dt=1
M27 23 19 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=11740 $dt=1
M28 45 43 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=2220 $dt=1
M29 38 36 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=4420 $dt=1
M30 31 29 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=9540 $dt=1
M31 24 22 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=11740 $dt=1
M32 83 43 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=1980 $dt=1
M33 81 36 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=4180 $dt=1
M34 79 29 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=9300 $dt=1
M35 77 22 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=11500 $dt=1
M36 12 44 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=2040 $dt=1
M37 13 37 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=4120 $dt=1
M38 14 30 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=9360 $dt=1
M39 15 23 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=11440 $dt=1
M40 12 45 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=2040 $dt=1
M41 13 38 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=4120 $dt=1
M42 14 31 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=9360 $dt=1
M43 15 24 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=11440 $dt=1
M44 83 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=2040 $dt=1
M45 81 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=4120 $dt=1
M46 79 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=9360 $dt=1
M47 77 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=11440 $dt=1
M48 46 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=2010 $dt=1
M49 39 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=4150 $dt=1
M50 32 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=9330 $dt=1
M51 25 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=11470 $dt=1
M52 5 43 46 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=2010 $dt=1
M53 5 36 39 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=4150 $dt=1
M54 5 29 32 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=9330 $dt=1
M55 5 22 25 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=11470 $dt=1
M56 47 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=2230 $dt=1
M57 40 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=4410 $dt=1
M58 33 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=9550 $dt=1
M59 26 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=11730 $dt=1
M60 5 1 47 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=2230 $dt=1
M61 5 2 40 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=4410 $dt=1
M62 5 3 33 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=9550 $dt=1
M63 5 4 26 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=11730 $dt=1
M64 18 46 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=2230 $dt=1
M65 17 39 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=4410 $dt=1
M66 19 32 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=9550 $dt=1
M67 16 25 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=11730 $dt=1
M68 5 47 18 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=2230 $dt=1
M69 5 40 17 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=4410 $dt=1
M70 5 33 19 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=9550 $dt=1
M71 5 26 16 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=11730 $dt=1
.ends FA_4bit

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small 1 2 3 4
** N=4 EP=4 FDC=2
X0 1 M1_PO_CDNS_16 $T=950 1780 0 90 $X=830 $Y=1680
X1 2 3 cellTmpl_CDNS_18 $T=120 140 0 0 $X=0 $Y=0
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7353 scb=0.0117274 scc=0.000445561 $X=1070 $Y=980 $dt=0
M1 4 1 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8675 scb=0.0146094 scc=0.000688105 $X=1070 $Y=2220 $dt=1
.ends INV_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 10badder                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 10badder 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 64
+ 65 66 67 68 69 70 149 150 151 152
+ 153 154 155 256 257 266 267
*.DEVICECLIMB
** N=267 EP=77 FDC=483
X0 2 M3_M2_CDNS_1 $T=52330 32180 0 90 $X=52080 $Y=32100
X1 35 M3_M2_CDNS_1 $T=52330 46820 0 90 $X=52080 $Y=46740
X2 36 M3_M2_CDNS_1 $T=53480 29020 0 0 $X=53400 $Y=28770
X3 37 M3_M2_CDNS_1 $T=53480 43660 0 0 $X=53400 $Y=43410
X4 38 M3_M2_CDNS_1 $T=54270 29810 0 90 $X=54020 $Y=29730
X5 39 M3_M2_CDNS_1 $T=54270 44450 0 90 $X=54020 $Y=44370
X6 36 M3_M2_CDNS_1 $T=55540 26280 0 0 $X=55460 $Y=26030
X7 37 M3_M2_CDNS_1 $T=55540 40920 0 0 $X=55460 $Y=40670
X8 40 M3_M2_CDNS_1 $T=55730 21200 0 90 $X=55480 $Y=21120
X9 41 M3_M2_CDNS_1 $T=55730 35840 0 90 $X=55480 $Y=35760
X10 42 M3_M2_CDNS_1 $T=56210 23810 0 90 $X=55960 $Y=23730
X11 43 M3_M2_CDNS_1 $T=56210 38450 0 90 $X=55960 $Y=38370
X12 44 M3_M2_CDNS_1 $T=56050 31070 0 0 $X=55970 $Y=30820
X13 45 M3_M2_CDNS_1 $T=56050 45710 0 0 $X=55970 $Y=45460
X14 46 M3_M2_CDNS_1 $T=56240 34220 0 0 $X=56160 $Y=33970
X15 47 M3_M2_CDNS_1 $T=56240 48860 0 0 $X=56160 $Y=48610
X16 13 M3_M2_CDNS_1 $T=57660 26200 0 90 $X=57410 $Y=26120
X17 11 M3_M2_CDNS_1 $T=57660 33520 0 90 $X=57410 $Y=33440
X18 10 M3_M2_CDNS_1 $T=57660 40840 0 90 $X=57410 $Y=40760
X19 8 M3_M2_CDNS_1 $T=57660 48160 0 90 $X=57410 $Y=48080
X20 7 M3_M2_CDNS_1 $T=57670 22770 0 90 $X=57420 $Y=22690
X21 12 M3_M2_CDNS_1 $T=57670 30070 0 90 $X=57420 $Y=29990
X22 6 M3_M2_CDNS_1 $T=57670 37410 0 90 $X=57420 $Y=37330
X23 9 M3_M2_CDNS_1 $T=57670 44710 0 90 $X=57420 $Y=44630
X24 44 M3_M2_CDNS_1 $T=62950 31240 0 90 $X=62700 $Y=31160
X25 45 M3_M2_CDNS_1 $T=62950 45880 0 90 $X=62700 $Y=45800
X26 42 M3_M2_CDNS_1 $T=63400 23460 0 0 $X=63320 $Y=23210
X27 43 M3_M2_CDNS_1 $T=63400 38100 0 0 $X=63320 $Y=37850
X28 40 M3_M2_CDNS_1 $T=63720 21760 0 0 $X=63640 $Y=21510
X29 41 M3_M2_CDNS_1 $T=63720 36400 0 0 $X=63640 $Y=36150
X30 38 M3_M2_CDNS_1 $T=63820 29420 0 0 $X=63740 $Y=29170
X31 39 M3_M2_CDNS_1 $T=63820 44060 0 0 $X=63740 $Y=43810
X32 36 M2_M1_CDNS_2 $T=53480 29020 0 0 $X=53400 $Y=28770
X33 37 M2_M1_CDNS_2 $T=53480 43660 0 0 $X=53400 $Y=43410
X34 46 M2_M1_CDNS_2 $T=56240 34220 0 0 $X=56160 $Y=33970
X35 47 M2_M1_CDNS_2 $T=56240 48860 0 0 $X=56160 $Y=48610
X36 44 M2_M1_CDNS_2 $T=62950 31240 0 90 $X=62700 $Y=31160
X37 45 M2_M1_CDNS_2 $T=62950 45880 0 90 $X=62700 $Y=45800
X38 42 M2_M1_CDNS_2 $T=63400 23460 0 0 $X=63320 $Y=23210
X39 43 M2_M1_CDNS_2 $T=63400 38100 0 0 $X=63320 $Y=37850
X40 40 M2_M1_CDNS_2 $T=63720 21760 0 0 $X=63640 $Y=21510
X41 41 M2_M1_CDNS_2 $T=63720 36400 0 0 $X=63640 $Y=36150
X42 38 M2_M1_CDNS_2 $T=63820 29420 0 0 $X=63740 $Y=29170
X43 39 M2_M1_CDNS_2 $T=63820 44060 0 0 $X=63740 $Y=43810
X44 35 M4_M3_CDNS_6 $T=51080 34160 0 0 $X=51000 $Y=33910
X45 48 M4_M3_CDNS_6 $T=56340 32800 0 0 $X=56260 $Y=32550
X46 49 M4_M3_CDNS_6 $T=56340 47440 0 0 $X=56260 $Y=47190
X47 50 M4_M3_CDNS_6 $T=57240 50840 0 0 $X=57160 $Y=50590
X48 51 M4_M3_CDNS_6 $T=72650 52420 0 90 $X=72400 $Y=52340
X49 35 M4_M3_CDNS_6 $T=78550 36430 0 0 $X=78470 $Y=36180
X50 51 M4_M3_CDNS_6 $T=79400 52420 0 90 $X=79150 $Y=52340
X51 48 M4_M3_CDNS_6 $T=86760 34460 0 0 $X=86680 $Y=34210
X52 49 M4_M3_CDNS_6 $T=86760 49100 0 0 $X=86680 $Y=48850
X53 35 M4_M3_CDNS_8 $T=51140 36930 0 0 $X=51060 $Y=36800
X54 35 M3_M2_CDNS_9 $T=51080 34160 0 0 $X=51000 $Y=33910
X55 48 M3_M2_CDNS_9 $T=56340 32800 0 0 $X=56260 $Y=32550
X56 49 M3_M2_CDNS_9 $T=56340 47440 0 0 $X=56260 $Y=47190
X57 50 M3_M2_CDNS_9 $T=57240 50840 0 0 $X=57160 $Y=50590
X58 51 M3_M2_CDNS_9 $T=72650 52420 0 90 $X=72400 $Y=52340
X59 35 M3_M2_CDNS_9 $T=78550 36430 0 0 $X=78470 $Y=36180
X60 51 M3_M2_CDNS_9 $T=79400 52420 0 90 $X=79150 $Y=52340
X61 48 M3_M2_CDNS_9 $T=86760 34460 0 0 $X=86680 $Y=34210
X62 49 M3_M2_CDNS_9 $T=86760 49100 0 0 $X=86680 $Y=48850
X63 35 M2_M1_CDNS_10 $T=51080 34160 0 0 $X=51000 $Y=33910
X64 2 M2_M1_CDNS_10 $T=52330 32180 0 90 $X=52080 $Y=32100
X65 35 M2_M1_CDNS_10 $T=52330 46820 0 90 $X=52080 $Y=46740
X66 38 M2_M1_CDNS_10 $T=54270 29810 0 90 $X=54020 $Y=29730
X67 39 M2_M1_CDNS_10 $T=54270 44450 0 90 $X=54020 $Y=44370
X68 36 M2_M1_CDNS_10 $T=55540 26280 0 0 $X=55460 $Y=26030
X69 37 M2_M1_CDNS_10 $T=55540 40920 0 0 $X=55460 $Y=40670
X70 40 M2_M1_CDNS_10 $T=55730 21200 0 90 $X=55480 $Y=21120
X71 41 M2_M1_CDNS_10 $T=55730 35840 0 90 $X=55480 $Y=35760
X72 42 M2_M1_CDNS_10 $T=56210 23810 0 90 $X=55960 $Y=23730
X73 43 M2_M1_CDNS_10 $T=56210 38450 0 90 $X=55960 $Y=38370
X74 44 M2_M1_CDNS_10 $T=56050 31070 0 0 $X=55970 $Y=30820
X75 45 M2_M1_CDNS_10 $T=56050 45710 0 0 $X=55970 $Y=45460
X76 48 M2_M1_CDNS_10 $T=56340 32800 0 0 $X=56260 $Y=32550
X77 49 M2_M1_CDNS_10 $T=56340 47440 0 0 $X=56260 $Y=47190
X78 50 M2_M1_CDNS_10 $T=57240 50840 0 0 $X=57160 $Y=50590
X79 13 M2_M1_CDNS_10 $T=57660 26200 0 90 $X=57410 $Y=26120
X80 11 M2_M1_CDNS_10 $T=57660 33520 0 90 $X=57410 $Y=33440
X81 10 M2_M1_CDNS_10 $T=57660 40840 0 90 $X=57410 $Y=40760
X82 8 M2_M1_CDNS_10 $T=57660 48160 0 90 $X=57410 $Y=48080
X83 7 M2_M1_CDNS_10 $T=57670 22770 0 90 $X=57420 $Y=22690
X84 12 M2_M1_CDNS_10 $T=57670 30070 0 90 $X=57420 $Y=29990
X85 6 M2_M1_CDNS_10 $T=57670 37410 0 90 $X=57420 $Y=37330
X86 9 M2_M1_CDNS_10 $T=57670 44710 0 90 $X=57420 $Y=44630
X87 51 M2_M1_CDNS_10 $T=72650 52420 0 90 $X=72400 $Y=52340
X88 35 M2_M1_CDNS_10 $T=78550 36430 0 0 $X=78470 $Y=36180
X89 51 M2_M1_CDNS_10 $T=79400 52420 0 90 $X=79150 $Y=52340
X90 48 M2_M1_CDNS_10 $T=86760 34460 0 0 $X=86680 $Y=34210
X91 49 M2_M1_CDNS_10 $T=86760 49100 0 0 $X=86680 $Y=48850
X92 3 M2_M1_CDNS_11 $T=50480 50560 0 0 $X=50400 $Y=50430
X93 3 M2_M1_CDNS_11 $T=51590 45750 0 90 $X=51460 $Y=45670
X94 46 M2_M1_CDNS_11 $T=53210 27000 0 0 $X=53130 $Y=26870
X95 47 M2_M1_CDNS_11 $T=53210 41640 0 0 $X=53130 $Y=41510
X96 52 M2_M1_CDNS_11 $T=53230 23140 0 0 $X=53150 $Y=23010
X97 53 M2_M1_CDNS_11 $T=53230 37780 0 0 $X=53150 $Y=37650
X98 3 M2_M1_CDNS_11 $T=62920 24380 0 0 $X=62840 $Y=24250
X99 3 M2_M1_CDNS_11 $T=62920 39020 0 0 $X=62840 $Y=38890
X100 3 M2_M1_CDNS_11 $T=62930 31710 0 0 $X=62850 $Y=31580
X101 3 M2_M1_CDNS_11 $T=62930 46350 0 0 $X=62850 $Y=46220
X102 2 M1_PO_CDNS_13 $T=52330 32180 0 90 $X=52080 $Y=32080
X103 35 M1_PO_CDNS_13 $T=52330 46820 0 90 $X=52080 $Y=46720
X104 38 M1_PO_CDNS_13 $T=54270 29810 0 90 $X=54020 $Y=29710
X105 39 M1_PO_CDNS_13 $T=54270 44450 0 90 $X=54020 $Y=44350
X106 36 M1_PO_CDNS_13 $T=55540 26280 0 0 $X=55440 $Y=26030
X107 37 M1_PO_CDNS_13 $T=55540 40920 0 0 $X=55440 $Y=40670
X108 40 M1_PO_CDNS_13 $T=55730 21200 0 90 $X=55480 $Y=21100
X109 41 M1_PO_CDNS_13 $T=55730 35840 0 90 $X=55480 $Y=35740
X110 44 M1_PO_CDNS_13 $T=56050 31070 0 0 $X=55950 $Y=30820
X111 45 M1_PO_CDNS_13 $T=56050 45710 0 0 $X=55950 $Y=45460
X112 42 M1_PO_CDNS_13 $T=56210 23810 0 90 $X=55960 $Y=23710
X113 43 M1_PO_CDNS_13 $T=56210 38450 0 90 $X=55960 $Y=38350
X114 48 M1_PO_CDNS_13 $T=56340 32800 0 0 $X=56240 $Y=32550
X115 49 M1_PO_CDNS_13 $T=56340 47440 0 0 $X=56240 $Y=47190
X116 13 M1_PO_CDNS_13 $T=57660 26200 0 90 $X=57410 $Y=26100
X117 11 M1_PO_CDNS_13 $T=57660 33520 0 90 $X=57410 $Y=33420
X118 10 M1_PO_CDNS_13 $T=57660 40840 0 90 $X=57410 $Y=40740
X119 8 M1_PO_CDNS_13 $T=57660 48160 0 90 $X=57410 $Y=48060
X120 7 M1_PO_CDNS_13 $T=57670 22770 0 90 $X=57420 $Y=22670
X121 12 M1_PO_CDNS_13 $T=57670 30070 0 90 $X=57420 $Y=29970
X122 6 M1_PO_CDNS_13 $T=57670 37410 0 90 $X=57420 $Y=37310
X123 9 M1_PO_CDNS_13 $T=57670 44710 0 90 $X=57420 $Y=44610
X124 35 M1_PO_CDNS_13 $T=78550 36430 0 0 $X=78450 $Y=36180
X125 46 M3_M2_CDNS_14 $T=50730 34460 0 0 $X=50650 $Y=34330
X126 47 M3_M2_CDNS_14 $T=50800 49100 0 0 $X=50720 $Y=48970
X127 2 M3_M2_CDNS_14 $T=51610 22610 0 0 $X=51530 $Y=22480
X128 52 M1_PO_CDNS_15 $T=53520 24980 0 90 $X=53270 $Y=24880
X129 53 M1_PO_CDNS_15 $T=53520 39620 0 90 $X=53270 $Y=39520
X130 14 M1_PO_CDNS_15 $T=64110 23330 0 0 $X=64010 $Y=23080
X131 18 M1_PO_CDNS_15 $T=64110 37970 0 0 $X=64010 $Y=37720
X132 14 M1_PO_CDNS_15 $T=65950 23850 0 90 $X=65700 $Y=23750
X133 18 M1_PO_CDNS_15 $T=65950 38490 0 90 $X=65700 $Y=38390
X134 2 M1_PO_CDNS_15 $T=78510 22370 0 0 $X=78410 $Y=22120
X135 54 M1_PO_CDNS_16 $T=53270 31100 0 0 $X=53170 $Y=30980
X136 55 M1_PO_CDNS_16 $T=53270 45740 0 0 $X=53170 $Y=45620
X137 56 M1_PO_CDNS_16 $T=53550 23450 0 0 $X=53450 $Y=23330
X138 57 M1_PO_CDNS_16 $T=53550 38090 0 0 $X=53450 $Y=37970
X139 58 M1_PO_CDNS_16 $T=53840 25910 0 0 $X=53740 $Y=25790
X140 59 M1_PO_CDNS_16 $T=53840 40550 0 0 $X=53740 $Y=40430
X141 52 M2_M1_CDNS_17 $T=53520 24980 0 90 $X=53270 $Y=24900
X142 53 M2_M1_CDNS_17 $T=53520 39620 0 90 $X=53270 $Y=39540
X143 14 M2_M1_CDNS_17 $T=64110 23330 0 0 $X=64030 $Y=23080
X144 18 M2_M1_CDNS_17 $T=64110 37970 0 0 $X=64030 $Y=37720
X145 14 M2_M1_CDNS_17 $T=65950 23850 0 90 $X=65700 $Y=23770
X146 18 M2_M1_CDNS_17 $T=65950 38490 0 90 $X=65700 $Y=38410
X147 2 M2_M1_CDNS_17 $T=78510 22370 0 0 $X=78430 $Y=22120
X148 3 4 40 56 42 172 NAND_1X_small $T=53960 20720 0 0 $X=53530 $Y=20700
X149 3 4 36 58 52 171 NAND_1X_small $T=55940 28040 0 180 $X=53530 $Y=24260
X150 3 4 38 54 44 170 NAND_1X_small $T=53960 28040 0 0 $X=53530 $Y=28020
X151 3 4 41 57 43 169 NAND_1X_small $T=53960 35360 0 0 $X=53530 $Y=35340
X152 3 4 37 59 53 168 NAND_1X_small $T=55940 42680 0 180 $X=53530 $Y=38900
X153 3 4 39 55 45 167 NAND_1X_small $T=53960 42680 0 0 $X=53530 $Y=42660
X154 3 4 14 7 42 85 86 187 265 188 XOR1 $T=56070 20720 0 0 $X=56130 $Y=20700
X155 3 4 15 13 40 83 84 185 264 186 XOR1 $T=56070 28040 1 0 $X=56130 $Y=24260
X156 3 4 16 12 44 81 82 183 263 184 XOR1 $T=56070 28040 0 0 $X=56130 $Y=28020
X157 3 4 17 11 38 79 80 181 262 182 XOR1 $T=56070 35360 1 0 $X=56130 $Y=31580
X158 3 4 18 6 43 77 78 179 261 180 XOR1 $T=56070 35360 0 0 $X=56130 $Y=35340
X159 3 4 19 10 41 75 76 177 260 178 XOR1 $T=56070 42680 1 0 $X=56130 $Y=38900
X160 3 4 20 9 45 73 74 175 259 176 XOR1 $T=56070 42680 0 0 $X=56130 $Y=42660
X161 3 4 21 8 39 71 72 173 258 174 XOR1 $T=56070 50000 1 0 $X=56130 $Y=46220
X162 5 3 1 4 50 22 51 66 69 70
+ 64 65 67 68 256 257 full_adder1_small $T=50650 49970 0 0 $X=50670 $Y=49980
X163 24 3 23 4 51 33 34 151 154 155
+ 149 150 152 153 266 267 full_adder1_small $T=72610 49970 0 0 $X=72630 $Y=49980
X164 46 48 3 4 2 35 62 63 158 159
+ 254 255 MUX_2to1___2X $T=56190 30160 0 180 $X=50640 $Y=31580
X165 47 49 3 4 35 50 60 61 156 157
+ 252 253 MUX_2to1___2X $T=56190 44800 0 180 $X=50640 $Y=46220
X166 14 13 12 11 3 7 4 15 16 17
+ 2 25 28 27 26 48 140 138 139 FA_4bit $T=64900 20820 0 0 $X=64250 $Y=20700
X167 18 10 9 8 3 6 4 19 20 21
+ 35 32 31 30 29 49 109 107 108 FA_4bit $T=64900 35460 0 0 $X=64250 $Y=35340
X168 56 3 4 52 INV_1X_small $T=51530 20700 0 0 $X=51530 $Y=20700
X169 58 3 4 46 INV_1X_small $T=51530 28060 1 0 $X=51530 $Y=24260
X170 54 3 4 36 INV_1X_small $T=51530 28020 0 0 $X=51530 $Y=28020
X171 57 3 4 53 INV_1X_small $T=51530 35340 0 0 $X=51530 $Y=35340
X172 59 3 4 47 INV_1X_small $T=51530 42700 1 0 $X=51530 $Y=38900
X173 55 3 4 37 INV_1X_small $T=51530 42660 0 0 $X=51530 $Y=42660
M0 64 5 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6612 scb=0.0167915 scc=0.000377457 $X=51440 $Y=52320 $dt=1
M1 58 52 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=25230 $dt=1
M2 59 53 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=39870 $dt=1
M3 56 40 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=23050 $dt=1
M4 54 38 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=30370 $dt=1
M5 57 41 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=37690 $dt=1
M6 55 39 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=45010 $dt=1
M7 3 36 58 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=25230 $dt=1
M8 3 37 59 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=39870 $dt=1
M9 3 42 56 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=23050 $dt=1
M10 3 44 54 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=30370 $dt=1
M11 3 43 57 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=37690 $dt=1
M12 3 45 55 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=45010 $dt=1
M13 85 14 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=23040 $dt=1
M14 83 15 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=25240 $dt=1
M15 81 16 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=30360 $dt=1
M16 79 17 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=32560 $dt=1
M17 77 18 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=37680 $dt=1
M18 75 19 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=39880 $dt=1
M19 73 20 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=45000 $dt=1
M20 71 21 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=47200 $dt=1
M21 86 7 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=23040 $dt=1
M22 84 13 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=25240 $dt=1
M23 82 12 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=30360 $dt=1
M24 80 11 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=32560 $dt=1
M25 78 6 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=37680 $dt=1
M26 76 10 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=39880 $dt=1
M27 74 9 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=45000 $dt=1
M28 72 8 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=47200 $dt=1
M29 265 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=22800 $dt=1
M30 264 13 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=25000 $dt=1
M31 263 12 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=30120 $dt=1
M32 262 11 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=32320 $dt=1
M33 261 6 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=37440 $dt=1
M34 260 10 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=39640 $dt=1
M35 259 9 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=44760 $dt=1
M36 258 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=46960 $dt=1
M37 42 85 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=22860 $dt=1
M38 40 83 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=24940 $dt=1
M39 44 81 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=30180 $dt=1
M40 38 79 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=32260 $dt=1
M41 43 77 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=37500 $dt=1
M42 41 75 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=39580 $dt=1
M43 45 73 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=44820 $dt=1
M44 39 71 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=46900 $dt=1
M45 42 86 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=22860 $dt=1
M46 40 84 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=24940 $dt=1
M47 44 82 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=30180 $dt=1
M48 38 80 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=32260 $dt=1
M49 43 78 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=37500 $dt=1
M50 41 76 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=39580 $dt=1
M51 45 74 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=44820 $dt=1
M52 39 72 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=46900 $dt=1
M53 265 14 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=22860 $dt=1
M54 264 15 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=24940 $dt=1
M55 263 16 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=30180 $dt=1
M56 262 17 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=32260 $dt=1
M57 261 18 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=37500 $dt=1
M58 260 19 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=39580 $dt=1
M59 259 20 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=44820 $dt=1
M60 258 21 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=46900 $dt=1
M61 34 154 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=93310 $Y=52330 $dt=1
M62 3 155 34 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=93720 $Y=52330 $dt=1
.ends 10badder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_46                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_46 1 2 3 5
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=660 $Y=760 $dt=0
.ends cellTmpl_CDNS_46

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 1 M1_PO_CDNS_16 $T=700 2040 0 90 $X=580 $Y=1940
X1 2 3 1 4 cellTmpl_CDNS_46 $T=120 140 0 0 $X=0 $Y=0
.ends INV_1X_small_layout

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_16 $T=640 1830 0 90 $X=520 $Y=1730
X1 6 M1_PO_CDNS_16 $T=1940 640 0 0 $X=1840 $Y=520
X2 3 1 6 3 nmos1v_CDNS_19 $T=710 860 0 0 $X=290 $Y=660
X3 4 6 5 3 nmos1v_CDNS_19 $T=1890 860 0 0 $X=1470 $Y=660
X4 2 3 cellTmpl_CDNS_21 $T=120 140 0 0 $X=0 $Y=0
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=710 $Y=860 $dt=0
M1 5 6 4 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1890 $Y=860 $dt=0
.ends ph1p3_clk_part

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_48                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_48 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_48

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_MSDFF                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_MSDFF 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17
*.DEVICECLIMB
** N=18 EP=17 FDC=15
X0 7 M3_M2_CDNS_1 $T=1140 2170 0 90 $X=890 $Y=2090
X1 8 M3_M2_CDNS_1 $T=3910 970 0 0 $X=3830 $Y=720
X2 9 M3_M2_CDNS_1 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X3 7 M3_M2_CDNS_1 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X4 7 M3_M2_CDNS_1 $T=8100 2170 0 90 $X=7850 $Y=2090
X5 9 M3_M2_CDNS_1 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X6 8 M3_M2_CDNS_1 $T=9760 1890 0 0 $X=9680 $Y=1640
X7 7 M2_M1_CDNS_2 $T=1140 2170 0 90 $X=890 $Y=2090
X8 8 M2_M1_CDNS_2 $T=3910 970 0 0 $X=3830 $Y=720
X9 9 M2_M1_CDNS_2 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X10 7 M2_M1_CDNS_2 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X11 9 M2_M1_CDNS_2 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X12 8 M2_M1_CDNS_2 $T=9760 1890 0 0 $X=9680 $Y=1640
X13 1 M4_M3_CDNS_6 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X14 1 M4_M3_CDNS_6 $T=5110 3310 0 0 $X=5030 $Y=3060
X15 1 M3_M2_CDNS_9 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X16 1 M3_M2_CDNS_9 $T=5110 3310 0 0 $X=5030 $Y=3060
X17 1 M2_M1_CDNS_10 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X18 1 M2_M1_CDNS_10 $T=5110 3310 0 0 $X=5030 $Y=3060
X19 7 M2_M1_CDNS_10 $T=8100 2170 0 90 $X=7850 $Y=2090
X20 2 M2_M1_CDNS_11 $T=430 2010 0 0 $X=350 $Y=1880
X21 10 M2_M1_CDNS_11 $T=1110 -1470 0 0 $X=1030 $Y=-1600
X22 2 M2_M1_CDNS_11 $T=2790 -1820 0 0 $X=2710 $Y=-1950
X23 11 M2_M1_CDNS_11 $T=4150 -1460 0 0 $X=4070 $Y=-1590
X24 6 M2_M1_CDNS_11 $T=5200 -2030 0 0 $X=5120 $Y=-2160
X25 10 M2_M1_CDNS_11 $T=5310 1560 0 90 $X=5180 $Y=1480
X26 11 M2_M1_CDNS_11 $T=5670 -1460 0 90 $X=5540 $Y=-1540
X27 12 M2_M1_CDNS_11 $T=6280 1490 0 0 $X=6200 $Y=1360
X28 13 M2_M1_CDNS_11 $T=7300 1510 0 90 $X=7170 $Y=1430
X29 12 M2_M1_CDNS_11 $T=7850 -2080 0 0 $X=7770 $Y=-2210
X30 13 M2_M1_CDNS_11 $T=9400 1510 0 90 $X=9270 $Y=1430
X31 6 M2_M1_CDNS_11 $T=9770 -2060 0 0 $X=9690 $Y=-2190
X32 7 M1_PO_CDNS_13 $T=8100 2170 0 90 $X=7850 $Y=2070
X33 8 1 3 10 12 18 NAND2_1X_small $T=3680 -70 0 0 $X=3800 $Y=0
X34 4 1 3 10 INV_1X_small_layout $T=0 40 1 0 $X=0 $Y=-3760
X35 2 1 3 7 INV_1X_small_layout $T=0 0 0 0 $X=0 $Y=0
X36 6 1 3 11 INV_1X_small_layout $T=4800 40 1 0 $X=4800 $Y=-3760
X37 12 1 3 13 INV_1X_small_layout $T=6200 0 0 0 $X=6200 $Y=0
X38 9 1 3 6 INV_1X_small_layout $T=8600 40 1 0 $X=8600 $Y=-3760
X39 2 1 3 5 8 14 ph1p3_clk_part $T=1400 0 0 0 $X=1400 $Y=0
X40 2 1 3 11 9 15 ph1p3_clk_part $T=2400 40 1 0 $X=2400 $Y=-3760
X41 7 1 3 12 9 16 ph1p3_clk_part $T=6200 40 1 0 $X=6200 $Y=-3760
X42 7 1 3 13 8 17 ph1p3_clk_part $T=7600 0 0 0 $X=7600 $Y=0
X43 1 3 cellTmpl_CDNS_48 $T=1520 -100 1 0 $X=1400 $Y=-3760
.ends ph1p3_MSDFF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_49                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_49 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_49

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X_ph2p2                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X_ph2p2 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=12 EP=12 FDC=6
X0 7 M3_M2_CDNS_1 $T=430 2220 0 0 $X=350 $Y=1970
X1 7 M3_M2_CDNS_1 $T=1140 3180 0 0 $X=1060 $Y=2930
X2 7 M3_M2_CDNS_1 $T=2800 2490 0 0 $X=2720 $Y=2240
X3 7 M2_M1_CDNS_2 $T=1140 3180 0 0 $X=1060 $Y=2930
X4 7 M2_M1_CDNS_10 $T=430 2220 0 0 $X=350 $Y=1970
X5 7 M2_M1_CDNS_10 $T=2800 2490 0 0 $X=2720 $Y=2240
X6 7 M1_PO_CDNS_13 $T=430 2220 0 0 $X=330 $Y=1970
X7 7 M1_PO_CDNS_13 $T=2800 2490 0 0 $X=2700 $Y=2240
X8 1 M1_PO_CDNS_15 $T=1480 1720 0 0 $X=1380 $Y=1470
X9 1 M1_PO_CDNS_15 $T=2840 980 0 0 $X=2740 $Y=730
X10 1 M1_PO_CDNS_16 $T=860 1670 0 0 $X=760 $Y=1550
X11 2 M1_PO_CDNS_16 $T=1480 3130 0 0 $X=1380 $Y=3010
X12 5 M1_PO_CDNS_16 $T=4220 2040 0 0 $X=4120 $Y=1920
X13 8 M1_PO_CDNS_16 $T=4480 1550 0 90 $X=4360 $Y=1450
X14 1 M2_M1_CDNS_17 $T=1480 1720 0 0 $X=1400 $Y=1470
X15 1 M2_M1_CDNS_17 $T=2840 980 0 0 $X=2760 $Y=730
X16 4 7 9 4 nmos1v_CDNS_31 $T=2170 800 0 0 $X=1970 $Y=600
X17 8 5 10 4 nmos1v_CDNS_31 $T=3550 790 0 0 $X=3350 $Y=590
X18 8 2 9 4 nmos1v_CDNS_32 $T=1960 800 0 0 $X=1540 $Y=600
X19 4 1 10 4 nmos1v_CDNS_32 $T=3340 790 0 0 $X=2920 $Y=590
X20 3 4 1 7 8 6 cellTmpl_CDNS_43 $T=120 140 0 0 $X=0 $Y=0
X21 3 1 11 4 3 pmos1v_CDNS_44 $T=2170 2100 0 0 $X=1970 $Y=1900
X22 8 5 12 4 3 pmos1v_CDNS_44 $T=3550 2030 0 0 $X=3350 $Y=1830
X23 8 2 11 4 3 pmos1v_CDNS_45 $T=1960 2100 0 0 $X=1540 $Y=1900
X24 3 7 12 4 3 pmos1v_CDNS_45 $T=3340 2030 0 0 $X=2920 $Y=1830
M0 9 2 8 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1960 $Y=800 $dt=0
M1 4 7 9 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=2170 $Y=800 $dt=0
M2 10 1 4 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3340 $Y=790 $dt=0
M3 8 5 10 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3550 $Y=790 $dt=0
.ends MUX_2to1___2X_ph2p2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p2_processing_element                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p2_processing_element 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 77 78 79 81 83
+ 108 113 130 139 140 141 158 159 176 185
+ 190 191 194 211 212 213 330 332 333 334
+ 336 338 348 350 351 352 354 356 366 368
+ 369 370 372 374 505 691 697 703 760 761
+ 762 763
*.DEVICECLIMB
** N=789 EP=122 FDC=1597
X0 6 M3_M2_CDNS_1 $T=1860 60810 0 0 $X=1780 $Y=60560
X1 6 M3_M2_CDNS_1 $T=1870 68120 0 0 $X=1790 $Y=67870
X2 6 M3_M2_CDNS_1 $T=12100 60800 0 0 $X=12020 $Y=60550
X3 6 M3_M2_CDNS_1 $T=12100 68120 0 0 $X=12020 $Y=67870
X4 6 M3_M2_CDNS_1 $T=22340 68120 0 0 $X=22260 $Y=67870
X5 6 M3_M2_CDNS_1 $T=22350 60800 0 0 $X=22270 $Y=60550
X6 46 M3_M2_CDNS_1 $T=22980 34240 0 0 $X=22900 $Y=33990
X7 47 M3_M2_CDNS_1 $T=28400 24370 0 0 $X=28320 $Y=24120
X8 48 M3_M2_CDNS_1 $T=32190 56290 0 0 $X=32110 $Y=56040
X9 6 M3_M2_CDNS_1 $T=32580 60800 0 0 $X=32500 $Y=60550
X10 6 M3_M2_CDNS_1 $T=32580 68120 0 0 $X=32500 $Y=67870
X11 6 M3_M2_CDNS_1 $T=40360 10220 0 90 $X=40110 $Y=10140
X12 6 M3_M2_CDNS_1 $T=40340 24940 0 0 $X=40260 $Y=24690
X13 6 M3_M2_CDNS_1 $T=40370 17590 0 0 $X=40290 $Y=17340
X14 49 M3_M2_CDNS_1 $T=45710 34580 0 0 $X=45630 $Y=34330
X15 6 M3_M2_CDNS_1 $T=47620 54480 0 90 $X=47370 $Y=54400
X16 6 M3_M2_CDNS_1 $T=47800 38230 0 90 $X=47550 $Y=38150
X17 6 M3_M2_CDNS_1 $T=47870 10240 0 0 $X=47790 $Y=9990
X18 6 M3_M2_CDNS_1 $T=48260 51950 0 90 $X=48010 $Y=51870
X19 6 M3_M2_CDNS_1 $T=48260 45130 0 0 $X=48180 $Y=44880
X20 6 M3_M2_CDNS_1 $T=48690 16910 0 0 $X=48610 $Y=16660
X21 6 M3_M2_CDNS_1 $T=48860 24230 0 0 $X=48780 $Y=23980
X22 50 M2_M1_CDNS_2 $T=14700 34240 0 0 $X=14620 $Y=33990
X23 46 M2_M1_CDNS_2 $T=22980 34240 0 0 $X=22900 $Y=33990
X24 47 M2_M1_CDNS_2 $T=28400 24370 0 0 $X=28320 $Y=24120
X25 48 M2_M1_CDNS_2 $T=32190 56290 0 0 $X=32110 $Y=56040
X26 51 M2_M1_CDNS_2 $T=38820 45300 0 0 $X=38740 $Y=45050
X27 49 M2_M1_CDNS_2 $T=45710 34580 0 0 $X=45630 $Y=34330
X28 52 M5_M4_CDNS_3 $T=31030 6520 0 0 $X=30950 $Y=6390
X29 53 M5_M4_CDNS_3 $T=33450 34810 0 0 $X=33370 $Y=34680
X30 53 M5_M4_CDNS_3 $T=34490 38940 0 0 $X=34410 $Y=38810
X31 53 M5_M4_CDNS_3 $T=35140 50450 0 0 $X=35060 $Y=50320
X32 54 M5_M4_CDNS_3 $T=35270 23970 0 0 $X=35190 $Y=23840
X33 53 M5_M4_CDNS_3 $T=35630 42220 0 0 $X=35550 $Y=42090
X34 52 M5_M4_CDNS_3 $T=35740 16590 0 0 $X=35660 $Y=16460
X35 55 M5_M4_CDNS_3 $T=36550 34300 0 0 $X=36470 $Y=34170
X36 47 M5_M4_CDNS_3 $T=36920 33010 0 0 $X=36840 $Y=32880
X37 56 M5_M4_CDNS_3 $T=37650 13930 0 0 $X=37570 $Y=13800
X38 57 M5_M4_CDNS_3 $T=37800 9740 0 0 $X=37720 $Y=9610
X39 58 M5_M4_CDNS_3 $T=38000 8190 0 0 $X=37920 $Y=8060
X40 59 M5_M4_CDNS_3 $T=38690 18860 0 90 $X=38560 $Y=18780
X41 60 M5_M4_CDNS_3 $T=38750 26290 0 90 $X=38620 $Y=26210
X42 59 M5_M4_CDNS_3 $T=40200 18860 0 90 $X=40070 $Y=18780
X43 58 M5_M4_CDNS_3 $T=40300 8620 0 90 $X=40170 $Y=8540
X44 61 M5_M4_CDNS_3 $T=48360 8140 0 0 $X=48280 $Y=8010
X45 61 M5_M4_CDNS_3 $T=50330 8160 0 0 $X=50250 $Y=8030
X46 47 M5_M4_CDNS_3 $T=50340 37430 0 0 $X=50260 $Y=37300
X47 62 M3_M2_CDNS_4 $T=15150 34320 0 0 $X=15070 $Y=34070
X48 63 M3_M2_CDNS_4 $T=30360 48950 0 0 $X=30280 $Y=48700
X49 51 M3_M2_CDNS_4 $T=30540 30290 0 90 $X=30290 $Y=30210
X50 64 M3_M2_CDNS_4 $T=30920 28440 0 90 $X=30670 $Y=28360
X51 64 M3_M2_CDNS_4 $T=30920 23090 0 0 $X=30840 $Y=22840
X52 51 M3_M2_CDNS_4 $T=30960 32190 0 0 $X=30880 $Y=31940
X53 65 M3_M2_CDNS_4 $T=34240 15510 0 0 $X=34160 $Y=15260
X54 60 M3_M2_CDNS_4 $T=36070 26280 0 0 $X=35990 $Y=26030
X55 51 M3_M2_CDNS_4 $T=36600 41550 0 0 $X=36520 $Y=41300
X56 54 M3_M2_CDNS_4 $T=37800 29000 0 0 $X=37720 $Y=28750
X57 66 M3_M2_CDNS_4 $T=40600 12040 0 0 $X=40520 $Y=11790
X58 61 M3_M2_CDNS_4 $T=41660 8130 0 0 $X=41580 $Y=7880
X59 58 M3_M2_CDNS_4 $T=43120 8620 0 0 $X=43040 $Y=8370
X60 7 M3_M2_CDNS_4 $T=45720 13840 0 0 $X=45640 $Y=13590
X61 7 M3_M2_CDNS_4 $T=47400 30300 0 0 $X=47320 $Y=30050
X62 47 M3_M2_CDNS_4 $T=50830 40760 0 90 $X=50580 $Y=40680
X63 25 M3_M2_CDNS_4 $T=58260 1650 0 0 $X=58180 $Y=1400
X64 1 M4_M3_CDNS_5 $T=1480 56760 0 0 $X=1400 $Y=56510
X65 4 M4_M3_CDNS_5 $T=2350 44590 0 90 $X=2100 $Y=44510
X66 3 M4_M3_CDNS_5 $T=3900 48300 0 90 $X=3650 $Y=48220
X67 2 M4_M3_CDNS_5 $T=3940 58210 0 90 $X=3690 $Y=58130
X68 1 M4_M3_CDNS_5 $T=4250 65060 0 0 $X=4170 $Y=64810
X69 2 M4_M3_CDNS_5 $T=4250 72470 0 0 $X=4170 $Y=72220
X70 10 M4_M3_CDNS_5 $T=6840 58120 0 90 $X=6590 $Y=58040
X71 14 M4_M3_CDNS_5 $T=11380 56560 0 90 $X=11130 $Y=56480
X72 14 M4_M3_CDNS_5 $T=14490 65150 0 0 $X=14410 $Y=64900
X73 10 M4_M3_CDNS_5 $T=14490 72480 0 0 $X=14410 $Y=72230
X74 13 M4_M3_CDNS_5 $T=20420 56560 0 90 $X=20170 $Y=56480
X75 13 M4_M3_CDNS_5 $T=24730 65150 0 0 $X=24650 $Y=64900
X76 3 M4_M3_CDNS_5 $T=24730 72470 0 0 $X=24650 $Y=72220
X77 67 M4_M3_CDNS_5 $T=27620 26990 0 0 $X=27540 $Y=26740
X78 15 M4_M3_CDNS_5 $T=29230 56560 0 90 $X=28980 $Y=56480
X79 68 M4_M3_CDNS_5 $T=32470 34080 0 90 $X=32220 $Y=34000
X80 52 M4_M3_CDNS_5 $T=33670 6150 0 90 $X=33420 $Y=6070
X81 15 M4_M3_CDNS_5 $T=34970 65150 0 0 $X=34890 $Y=64900
X82 4 M4_M3_CDNS_5 $T=34970 72470 0 0 $X=34890 $Y=72220
X83 53 M4_M3_CDNS_5 $T=35130 53970 0 0 $X=35050 $Y=53720
X84 56 M4_M3_CDNS_5 $T=38220 15840 0 0 $X=38140 $Y=15590
X85 52 M4_M3_CDNS_5 $T=38250 22590 0 0 $X=38170 $Y=22340
X86 69 M4_M3_CDNS_5 $T=38270 21170 0 0 $X=38190 $Y=20920
X87 58 M4_M3_CDNS_5 $T=47280 7640 0 90 $X=47030 $Y=7560
X88 56 M4_M3_CDNS_5 $T=47850 15290 0 0 $X=47770 $Y=15040
X89 52 M4_M3_CDNS_5 $T=47850 23870 0 0 $X=47770 $Y=23620
X90 6 M4_M3_CDNS_5 $T=47980 9490 0 0 $X=47900 $Y=9240
X91 6 M4_M3_CDNS_5 $T=48880 2280 0 0 $X=48800 $Y=2030
X92 7 M4_M3_CDNS_5 $T=50250 45640 0 90 $X=50000 $Y=45560
X93 58 M4_M3_CDNS_5 $T=59660 13790 0 0 $X=59580 $Y=13540
X94 56 M4_M3_CDNS_5 $T=59660 21120 0 0 $X=59580 $Y=20870
X95 52 M4_M3_CDNS_5 $T=59660 28470 0 0 $X=59580 $Y=28220
X96 5 M4_M3_CDNS_6 $T=1340 55390 0 0 $X=1260 $Y=55140
X97 5 M4_M3_CDNS_6 $T=3450 61970 0 0 $X=3370 $Y=61720
X98 5 M4_M3_CDNS_6 $T=9870 69280 0 0 $X=9790 $Y=69030
X99 50 M4_M3_CDNS_6 $T=14700 34240 0 0 $X=14620 $Y=33990
X100 62 M4_M3_CDNS_6 $T=15150 34320 0 0 $X=15070 $Y=34070
X101 70 M4_M3_CDNS_6 $T=28040 20980 0 0 $X=27960 $Y=20730
X102 63 M4_M3_CDNS_6 $T=30360 48950 0 0 $X=30280 $Y=48700
X103 51 M4_M3_CDNS_6 $T=30540 30290 0 90 $X=30290 $Y=30210
X104 64 M4_M3_CDNS_6 $T=30920 28440 0 90 $X=30670 $Y=28360
X105 64 M4_M3_CDNS_6 $T=30920 23090 0 0 $X=30840 $Y=22840
X106 51 M4_M3_CDNS_6 $T=30960 32190 0 0 $X=30880 $Y=31940
X107 65 M4_M3_CDNS_6 $T=34240 15510 0 0 $X=34160 $Y=15260
X108 60 M4_M3_CDNS_6 $T=36070 26280 0 0 $X=35990 $Y=26030
X109 51 M4_M3_CDNS_6 $T=36600 41550 0 0 $X=36520 $Y=41300
X110 49 M4_M3_CDNS_6 $T=37620 30320 0 0 $X=37540 $Y=30070
X111 54 M4_M3_CDNS_6 $T=37800 29000 0 0 $X=37720 $Y=28750
X112 51 M4_M3_CDNS_6 $T=38820 45300 0 0 $X=38740 $Y=45050
X113 66 M4_M3_CDNS_6 $T=40600 12040 0 0 $X=40520 $Y=11790
X114 66 M4_M3_CDNS_6 $T=40600 13810 0 0 $X=40520 $Y=13560
X115 61 M4_M3_CDNS_6 $T=41660 8130 0 0 $X=41580 $Y=7880
X116 58 M4_M3_CDNS_6 $T=43120 8620 0 0 $X=43040 $Y=8370
X117 7 M4_M3_CDNS_6 $T=45720 13840 0 0 $X=45640 $Y=13590
X118 7 M4_M3_CDNS_6 $T=46890 13630 0 0 $X=46810 $Y=13380
X119 7 M4_M3_CDNS_6 $T=46900 20740 0 0 $X=46820 $Y=20490
X120 7 M4_M3_CDNS_6 $T=46910 28080 0 0 $X=46830 $Y=27830
X121 5 M4_M3_CDNS_6 $T=49180 4060 0 0 $X=49100 $Y=3810
X122 5 M4_M3_CDNS_6 $T=49180 11470 0 0 $X=49100 $Y=11220
X123 5 M4_M3_CDNS_6 $T=49180 18800 0 0 $X=49100 $Y=18550
X124 5 M4_M3_CDNS_6 $T=49180 26120 0 0 $X=49100 $Y=25870
X125 5 M4_M3_CDNS_6 $T=49180 33430 0 0 $X=49100 $Y=33180
X126 5 M4_M3_CDNS_6 $T=49180 40820 0 0 $X=49100 $Y=40570
X127 5 M4_M3_CDNS_6 $T=49180 48070 0 0 $X=49100 $Y=47820
X128 5 M4_M3_CDNS_6 $T=49180 54710 0 0 $X=49100 $Y=54460
X129 47 M4_M3_CDNS_6 $T=50830 40760 0 90 $X=50580 $Y=40680
X130 25 M4_M3_CDNS_6 $T=58260 1650 0 0 $X=58180 $Y=1400
X131 25 M4_M3_CDNS_6 $T=58670 9650 0 90 $X=58420 $Y=9570
X132 25 M4_M3_CDNS_6 $T=58670 12550 0 90 $X=58420 $Y=12470
X133 25 M4_M3_CDNS_6 $T=58670 16970 0 90 $X=58420 $Y=16890
X134 25 M4_M3_CDNS_6 $T=58670 19870 0 90 $X=58420 $Y=19790
X135 25 M4_M3_CDNS_6 $T=58670 24290 0 90 $X=58420 $Y=24210
X136 25 M4_M3_CDNS_6 $T=58670 27190 0 90 $X=58420 $Y=27110
X137 25 M4_M3_CDNS_6 $T=58670 31610 0 90 $X=58420 $Y=31530
X138 25 M4_M3_CDNS_6 $T=58670 38930 0 90 $X=58420 $Y=38850
X139 25 M4_M3_CDNS_6 $T=58670 46250 0 90 $X=58420 $Y=46170
X140 25 M4_M3_CDNS_6 $T=58670 53570 0 90 $X=58420 $Y=53490
X141 1 M5_M4_CDNS_7 $T=1480 56760 0 0 $X=1400 $Y=56510
X142 4 M5_M4_CDNS_7 $T=2350 44590 0 90 $X=2100 $Y=44510
X143 3 M5_M4_CDNS_7 $T=3900 48300 0 90 $X=3650 $Y=48220
X144 2 M5_M4_CDNS_7 $T=3940 58210 0 90 $X=3690 $Y=58130
X145 1 M5_M4_CDNS_7 $T=4250 65060 0 0 $X=4170 $Y=64810
X146 2 M5_M4_CDNS_7 $T=4250 72470 0 0 $X=4170 $Y=72220
X147 10 M5_M4_CDNS_7 $T=6840 58120 0 90 $X=6590 $Y=58040
X148 14 M5_M4_CDNS_7 $T=11380 56560 0 90 $X=11130 $Y=56480
X149 14 M5_M4_CDNS_7 $T=14490 65150 0 0 $X=14410 $Y=64900
X150 10 M5_M4_CDNS_7 $T=14490 72480 0 0 $X=14410 $Y=72230
X151 13 M5_M4_CDNS_7 $T=20420 56560 0 90 $X=20170 $Y=56480
X152 13 M5_M4_CDNS_7 $T=24730 65150 0 0 $X=24650 $Y=64900
X153 3 M5_M4_CDNS_7 $T=24730 72470 0 0 $X=24650 $Y=72220
X154 67 M5_M4_CDNS_7 $T=27620 26990 0 0 $X=27540 $Y=26740
X155 15 M5_M4_CDNS_7 $T=29230 56560 0 90 $X=28980 $Y=56480
X156 67 M5_M4_CDNS_7 $T=32380 35710 0 90 $X=32130 $Y=35630
X157 68 M5_M4_CDNS_7 $T=32470 34080 0 90 $X=32220 $Y=34000
X158 68 M5_M4_CDNS_7 $T=33360 32510 0 90 $X=33110 $Y=32430
X159 52 M5_M4_CDNS_7 $T=33670 6150 0 90 $X=33420 $Y=6070
X160 55 M5_M4_CDNS_7 $T=33880 28620 0 0 $X=33800 $Y=28370
X161 53 M5_M4_CDNS_7 $T=34010 30140 0 0 $X=33930 $Y=29890
X162 54 M5_M4_CDNS_7 $T=34370 21060 0 0 $X=34290 $Y=20810
X163 15 M5_M4_CDNS_7 $T=34970 65150 0 0 $X=34890 $Y=64900
X164 4 M5_M4_CDNS_7 $T=34970 72470 0 0 $X=34890 $Y=72220
X165 53 M5_M4_CDNS_7 $T=35130 53970 0 0 $X=35050 $Y=53720
X166 69 M5_M4_CDNS_7 $T=36160 20250 0 0 $X=36080 $Y=20000
X167 71 M5_M4_CDNS_7 $T=36500 13950 0 0 $X=36420 $Y=13700
X168 72 M5_M4_CDNS_7 $T=37400 32460 0 0 $X=37320 $Y=32210
X169 65 M5_M4_CDNS_7 $T=37820 20120 0 0 $X=37740 $Y=19870
X170 56 M5_M4_CDNS_7 $T=38220 15840 0 0 $X=38140 $Y=15590
X171 52 M5_M4_CDNS_7 $T=38250 22590 0 0 $X=38170 $Y=22340
X172 69 M5_M4_CDNS_7 $T=38270 21170 0 0 $X=38190 $Y=20920
X173 71 M5_M4_CDNS_7 $T=40460 17040 0 90 $X=40210 $Y=16960
X174 65 M5_M4_CDNS_7 $T=40660 20120 0 90 $X=40410 $Y=20040
X175 57 M5_M4_CDNS_7 $T=40730 9730 0 90 $X=40480 $Y=9650
X176 60 M5_M4_CDNS_7 $T=40560 26320 0 0 $X=40480 $Y=26070
X177 72 M5_M4_CDNS_7 $T=42630 35130 0 90 $X=42380 $Y=35050
X178 58 M5_M4_CDNS_7 $T=47280 7640 0 90 $X=47030 $Y=7560
X179 56 M5_M4_CDNS_7 $T=47850 15290 0 0 $X=47770 $Y=15040
X180 52 M5_M4_CDNS_7 $T=47850 23870 0 0 $X=47770 $Y=23620
X181 7 M5_M4_CDNS_7 $T=47890 45870 0 0 $X=47810 $Y=45620
X182 6 M5_M4_CDNS_7 $T=47980 9490 0 0 $X=47900 $Y=9240
X183 6 M5_M4_CDNS_7 $T=48880 2280 0 0 $X=48800 $Y=2030
X184 7 M5_M4_CDNS_7 $T=50250 45640 0 90 $X=50000 $Y=45560
X185 58 M5_M4_CDNS_7 $T=59660 13790 0 0 $X=59580 $Y=13540
X186 56 M5_M4_CDNS_7 $T=59660 21120 0 0 $X=59580 $Y=20870
X187 52 M5_M4_CDNS_7 $T=59660 28470 0 0 $X=59580 $Y=28220
X188 50 M4_M3_CDNS_8 $T=13710 9140 0 0 $X=13630 $Y=9010
X189 50 M4_M3_CDNS_8 $T=13710 17480 0 0 $X=13630 $Y=17350
X190 50 M4_M3_CDNS_8 $T=13710 19960 0 0 $X=13630 $Y=19830
X191 62 M4_M3_CDNS_8 $T=14090 21060 0 0 $X=14010 $Y=20930
X192 48 M4_M3_CDNS_8 $T=24590 43490 0 0 $X=24510 $Y=43360
X193 63 M4_M3_CDNS_8 $T=28000 27530 0 0 $X=27920 $Y=27400
X194 48 M4_M3_CDNS_8 $T=28120 30940 0 0 $X=28040 $Y=30810
X195 56 M4_M3_CDNS_8 $T=30320 6550 0 0 $X=30240 $Y=6420
X196 52 M4_M3_CDNS_8 $T=31030 8560 0 90 $X=30900 $Y=8480
X197 57 M4_M3_CDNS_8 $T=34270 8400 0 0 $X=34190 $Y=8270
X198 49 M4_M3_CDNS_8 $T=34570 23190 0 0 $X=34490 $Y=23060
X199 52 M4_M3_CDNS_8 $T=34690 12200 0 0 $X=34610 $Y=12070
X200 47 M4_M3_CDNS_8 $T=36100 30140 0 0 $X=36020 $Y=30010
X201 55 M4_M3_CDNS_8 $T=36540 37650 0 90 $X=36410 $Y=37570
X202 65 M4_M3_CDNS_8 $T=37250 15560 0 0 $X=37170 $Y=15430
X203 70 M4_M3_CDNS_8 $T=37310 22870 0 0 $X=37230 $Y=22740
X204 73 M4_M3_CDNS_8 $T=37550 19040 0 0 $X=37470 $Y=18910
X205 73 M4_M3_CDNS_8 $T=37670 21700 0 0 $X=37590 $Y=21570
X206 59 M4_M3_CDNS_8 $T=38370 9550 0 0 $X=38290 $Y=9420
X207 59 M4_M3_CDNS_8 $T=40710 21060 0 0 $X=40630 $Y=20930
X208 58 M4_M3_CDNS_8 $T=41120 2720 0 0 $X=41040 $Y=2590
X209 7 M4_M3_CDNS_8 $T=47400 30300 0 0 $X=47320 $Y=30170
X210 6 M4_M3_CDNS_8 $T=48170 14160 0 0 $X=48090 $Y=14030
X211 6 M4_M3_CDNS_8 $T=48170 17210 0 0 $X=48090 $Y=17080
X212 61 M4_M3_CDNS_8 $T=50910 13780 0 0 $X=50830 $Y=13650
X213 5 M3_M2_CDNS_9 $T=1340 55390 0 0 $X=1260 $Y=55140
X214 1 M3_M2_CDNS_9 $T=1480 56760 0 0 $X=1400 $Y=56510
X215 4 M3_M2_CDNS_9 $T=2350 44590 0 90 $X=2100 $Y=44510
X216 5 M3_M2_CDNS_9 $T=3450 61970 0 0 $X=3370 $Y=61720
X217 3 M3_M2_CDNS_9 $T=3900 48300 0 90 $X=3650 $Y=48220
X218 2 M3_M2_CDNS_9 $T=3940 58210 0 90 $X=3690 $Y=58130
X219 1 M3_M2_CDNS_9 $T=4250 65060 0 0 $X=4170 $Y=64810
X220 2 M3_M2_CDNS_9 $T=4250 72470 0 0 $X=4170 $Y=72220
X221 10 M3_M2_CDNS_9 $T=6840 58120 0 90 $X=6590 $Y=58040
X222 5 M3_M2_CDNS_9 $T=9870 69280 0 0 $X=9790 $Y=69030
X223 14 M3_M2_CDNS_9 $T=11380 56560 0 90 $X=11130 $Y=56480
X224 14 M3_M2_CDNS_9 $T=14490 65150 0 0 $X=14410 $Y=64900
X225 10 M3_M2_CDNS_9 $T=14490 72480 0 0 $X=14410 $Y=72230
X226 50 M3_M2_CDNS_9 $T=14700 34240 0 0 $X=14620 $Y=33990
X227 13 M3_M2_CDNS_9 $T=20420 56560 0 90 $X=20170 $Y=56480
X228 13 M3_M2_CDNS_9 $T=24730 65150 0 0 $X=24650 $Y=64900
X229 3 M3_M2_CDNS_9 $T=24730 72470 0 0 $X=24650 $Y=72220
X230 67 M3_M2_CDNS_9 $T=27620 26990 0 0 $X=27540 $Y=26740
X231 70 M3_M2_CDNS_9 $T=28040 20980 0 0 $X=27960 $Y=20730
X232 15 M3_M2_CDNS_9 $T=29230 56560 0 90 $X=28980 $Y=56480
X233 68 M3_M2_CDNS_9 $T=32470 34080 0 90 $X=32220 $Y=34000
X234 52 M3_M2_CDNS_9 $T=33670 6150 0 90 $X=33420 $Y=6070
X235 15 M3_M2_CDNS_9 $T=34970 65150 0 0 $X=34890 $Y=64900
X236 4 M3_M2_CDNS_9 $T=34970 72470 0 0 $X=34890 $Y=72220
X237 53 M3_M2_CDNS_9 $T=35130 53970 0 0 $X=35050 $Y=53720
X238 49 M3_M2_CDNS_9 $T=37620 30320 0 0 $X=37540 $Y=30070
X239 56 M3_M2_CDNS_9 $T=38220 15840 0 0 $X=38140 $Y=15590
X240 52 M3_M2_CDNS_9 $T=38250 22590 0 0 $X=38170 $Y=22340
X241 69 M3_M2_CDNS_9 $T=38270 21170 0 0 $X=38190 $Y=20920
X242 51 M3_M2_CDNS_9 $T=38820 45300 0 0 $X=38740 $Y=45050
X243 66 M3_M2_CDNS_9 $T=40600 13810 0 0 $X=40520 $Y=13560
X244 59 M3_M2_CDNS_9 $T=40710 21060 0 0 $X=40630 $Y=20810
X245 7 M3_M2_CDNS_9 $T=46890 13630 0 0 $X=46810 $Y=13380
X246 7 M3_M2_CDNS_9 $T=46900 20740 0 0 $X=46820 $Y=20490
X247 7 M3_M2_CDNS_9 $T=46910 28080 0 0 $X=46830 $Y=27830
X248 58 M3_M2_CDNS_9 $T=47280 7640 0 90 $X=47030 $Y=7560
X249 56 M3_M2_CDNS_9 $T=47850 15290 0 0 $X=47770 $Y=15040
X250 52 M3_M2_CDNS_9 $T=47850 23870 0 0 $X=47770 $Y=23620
X251 6 M3_M2_CDNS_9 $T=47980 9490 0 0 $X=47900 $Y=9240
X252 6 M3_M2_CDNS_9 $T=48880 2280 0 0 $X=48800 $Y=2030
X253 5 M3_M2_CDNS_9 $T=49180 4060 0 0 $X=49100 $Y=3810
X254 5 M3_M2_CDNS_9 $T=49180 11470 0 0 $X=49100 $Y=11220
X255 5 M3_M2_CDNS_9 $T=49180 18800 0 0 $X=49100 $Y=18550
X256 5 M3_M2_CDNS_9 $T=49180 26120 0 0 $X=49100 $Y=25870
X257 5 M3_M2_CDNS_9 $T=49180 33430 0 0 $X=49100 $Y=33180
X258 5 M3_M2_CDNS_9 $T=49180 40820 0 0 $X=49100 $Y=40570
X259 5 M3_M2_CDNS_9 $T=49180 48070 0 0 $X=49100 $Y=47820
X260 5 M3_M2_CDNS_9 $T=49180 54710 0 0 $X=49100 $Y=54460
X261 7 M3_M2_CDNS_9 $T=50250 45640 0 90 $X=50000 $Y=45560
X262 61 M3_M2_CDNS_9 $T=50910 13780 0 0 $X=50830 $Y=13530
X263 25 M3_M2_CDNS_9 $T=58670 9650 0 90 $X=58420 $Y=9570
X264 25 M3_M2_CDNS_9 $T=58670 12550 0 90 $X=58420 $Y=12470
X265 25 M3_M2_CDNS_9 $T=58670 16970 0 90 $X=58420 $Y=16890
X266 25 M3_M2_CDNS_9 $T=58670 19870 0 90 $X=58420 $Y=19790
X267 25 M3_M2_CDNS_9 $T=58670 24290 0 90 $X=58420 $Y=24210
X268 25 M3_M2_CDNS_9 $T=58670 27190 0 90 $X=58420 $Y=27110
X269 25 M3_M2_CDNS_9 $T=58670 31610 0 90 $X=58420 $Y=31530
X270 25 M3_M2_CDNS_9 $T=58670 38930 0 90 $X=58420 $Y=38850
X271 25 M3_M2_CDNS_9 $T=58670 46250 0 90 $X=58420 $Y=46170
X272 25 M3_M2_CDNS_9 $T=58670 53570 0 90 $X=58420 $Y=53490
X273 58 M3_M2_CDNS_9 $T=59660 13790 0 0 $X=59580 $Y=13540
X274 56 M3_M2_CDNS_9 $T=59660 21120 0 0 $X=59580 $Y=20870
X275 52 M3_M2_CDNS_9 $T=59660 28470 0 0 $X=59580 $Y=28220
X276 5 M2_M1_CDNS_10 $T=1340 55390 0 0 $X=1260 $Y=55140
X277 1 M2_M1_CDNS_10 $T=1480 56760 0 0 $X=1400 $Y=56510
X278 6 M2_M1_CDNS_10 $T=1860 60810 0 0 $X=1780 $Y=60560
X279 6 M2_M1_CDNS_10 $T=1870 68120 0 0 $X=1790 $Y=67870
X280 4 M2_M1_CDNS_10 $T=2350 44590 0 90 $X=2100 $Y=44510
X281 5 M2_M1_CDNS_10 $T=3450 61970 0 0 $X=3370 $Y=61720
X282 3 M2_M1_CDNS_10 $T=3900 48300 0 90 $X=3650 $Y=48220
X283 2 M2_M1_CDNS_10 $T=3940 58210 0 90 $X=3690 $Y=58130
X284 1 M2_M1_CDNS_10 $T=4250 65060 0 0 $X=4170 $Y=64810
X285 2 M2_M1_CDNS_10 $T=4250 72470 0 0 $X=4170 $Y=72220
X286 10 M2_M1_CDNS_10 $T=6840 58120 0 90 $X=6590 $Y=58040
X287 5 M2_M1_CDNS_10 $T=9870 69280 0 0 $X=9790 $Y=69030
X288 14 M2_M1_CDNS_10 $T=11380 56560 0 90 $X=11130 $Y=56480
X289 6 M2_M1_CDNS_10 $T=12100 60800 0 0 $X=12020 $Y=60550
X290 6 M2_M1_CDNS_10 $T=12100 68120 0 0 $X=12020 $Y=67870
X291 14 M2_M1_CDNS_10 $T=14490 65150 0 0 $X=14410 $Y=64900
X292 10 M2_M1_CDNS_10 $T=14490 72480 0 0 $X=14410 $Y=72230
X293 13 M2_M1_CDNS_10 $T=20420 56560 0 90 $X=20170 $Y=56480
X294 6 M2_M1_CDNS_10 $T=22340 68120 0 0 $X=22260 $Y=67870
X295 6 M2_M1_CDNS_10 $T=22350 60800 0 0 $X=22270 $Y=60550
X296 13 M2_M1_CDNS_10 $T=24730 65150 0 0 $X=24650 $Y=64900
X297 3 M2_M1_CDNS_10 $T=24730 72470 0 0 $X=24650 $Y=72220
X298 67 M2_M1_CDNS_10 $T=27620 26990 0 0 $X=27540 $Y=26740
X299 70 M2_M1_CDNS_10 $T=28040 20980 0 0 $X=27960 $Y=20730
X300 15 M2_M1_CDNS_10 $T=29230 56560 0 90 $X=28980 $Y=56480
X301 6 M2_M1_CDNS_10 $T=32580 60800 0 0 $X=32500 $Y=60550
X302 6 M2_M1_CDNS_10 $T=32580 68120 0 0 $X=32500 $Y=67870
X303 52 M2_M1_CDNS_10 $T=33670 6150 0 90 $X=33420 $Y=6070
X304 15 M2_M1_CDNS_10 $T=34970 65150 0 0 $X=34890 $Y=64900
X305 4 M2_M1_CDNS_10 $T=34970 72470 0 0 $X=34890 $Y=72220
X306 49 M2_M1_CDNS_10 $T=37620 30320 0 0 $X=37540 $Y=30070
X307 6 M2_M1_CDNS_10 $T=40360 10220 0 90 $X=40110 $Y=10140
X308 6 M2_M1_CDNS_10 $T=40340 24940 0 0 $X=40260 $Y=24690
X309 6 M2_M1_CDNS_10 $T=40370 17590 0 0 $X=40290 $Y=17340
X310 66 M2_M1_CDNS_10 $T=40600 13810 0 0 $X=40520 $Y=13560
X311 59 M2_M1_CDNS_10 $T=40710 21060 0 0 $X=40630 $Y=20810
X312 7 M2_M1_CDNS_10 $T=46890 13630 0 0 $X=46810 $Y=13380
X313 7 M2_M1_CDNS_10 $T=46900 20740 0 0 $X=46820 $Y=20490
X314 7 M2_M1_CDNS_10 $T=46910 28080 0 0 $X=46830 $Y=27830
X315 6 M2_M1_CDNS_10 $T=47620 54480 0 90 $X=47370 $Y=54400
X316 6 M2_M1_CDNS_10 $T=47800 38230 0 90 $X=47550 $Y=38150
X317 6 M2_M1_CDNS_10 $T=47870 10240 0 0 $X=47790 $Y=9990
X318 6 M2_M1_CDNS_10 $T=47980 9490 0 0 $X=47900 $Y=9240
X319 6 M2_M1_CDNS_10 $T=48260 51950 0 90 $X=48010 $Y=51870
X320 6 M2_M1_CDNS_10 $T=48260 45130 0 0 $X=48180 $Y=44880
X321 6 M2_M1_CDNS_10 $T=48690 16910 0 0 $X=48610 $Y=16660
X322 6 M2_M1_CDNS_10 $T=48860 24230 0 0 $X=48780 $Y=23980
X323 6 M2_M1_CDNS_10 $T=48880 2280 0 0 $X=48800 $Y=2030
X324 5 M2_M1_CDNS_10 $T=49180 4060 0 0 $X=49100 $Y=3810
X325 5 M2_M1_CDNS_10 $T=49180 11470 0 0 $X=49100 $Y=11220
X326 5 M2_M1_CDNS_10 $T=49180 18800 0 0 $X=49100 $Y=18550
X327 5 M2_M1_CDNS_10 $T=49180 26120 0 0 $X=49100 $Y=25870
X328 5 M2_M1_CDNS_10 $T=49180 33430 0 0 $X=49100 $Y=33180
X329 5 M2_M1_CDNS_10 $T=49180 40820 0 0 $X=49100 $Y=40570
X330 5 M2_M1_CDNS_10 $T=49180 48070 0 0 $X=49100 $Y=47820
X331 5 M2_M1_CDNS_10 $T=49180 54710 0 0 $X=49100 $Y=54460
X332 61 M2_M1_CDNS_10 $T=50910 13780 0 0 $X=50830 $Y=13530
X333 25 M2_M1_CDNS_10 $T=58670 9650 0 90 $X=58420 $Y=9570
X334 25 M2_M1_CDNS_10 $T=58670 12550 0 90 $X=58420 $Y=12470
X335 25 M2_M1_CDNS_10 $T=58670 16970 0 90 $X=58420 $Y=16890
X336 25 M2_M1_CDNS_10 $T=58670 19870 0 90 $X=58420 $Y=19790
X337 25 M2_M1_CDNS_10 $T=58670 24290 0 90 $X=58420 $Y=24210
X338 25 M2_M1_CDNS_10 $T=58670 27190 0 90 $X=58420 $Y=27110
X339 25 M2_M1_CDNS_10 $T=58670 31610 0 90 $X=58420 $Y=31530
X340 25 M2_M1_CDNS_10 $T=58670 38930 0 90 $X=58420 $Y=38850
X341 25 M2_M1_CDNS_10 $T=58670 46250 0 90 $X=58420 $Y=46170
X342 25 M2_M1_CDNS_10 $T=58670 53570 0 90 $X=58420 $Y=53490
X343 58 M2_M1_CDNS_10 $T=59660 13790 0 0 $X=59580 $Y=13540
X344 56 M2_M1_CDNS_10 $T=59660 21120 0 0 $X=59580 $Y=20870
X345 52 M2_M1_CDNS_10 $T=59660 28470 0 0 $X=59580 $Y=28220
X346 59 M2_M1_CDNS_11 $T=13960 1790 0 90 $X=13830 $Y=1710
X347 62 M2_M1_CDNS_11 $T=26670 45180 0 0 $X=26590 $Y=45050
X348 72 M2_M1_CDNS_11 $T=27600 31220 0 0 $X=27520 $Y=31090
X349 73 M2_M1_CDNS_11 $T=28050 6240 0 0 $X=27970 $Y=6110
X350 65 M2_M1_CDNS_11 $T=28100 13310 0 0 $X=28020 $Y=13180
X351 61 M2_M1_CDNS_11 $T=28110 10050 0 0 $X=28030 $Y=9920
X352 60 M2_M1_CDNS_11 $T=28410 16430 0 90 $X=28280 $Y=16350
X353 68 M2_M1_CDNS_11 $T=35470 34490 0 0 $X=35390 $Y=34360
X354 66 M2_M1_CDNS_11 $T=35820 2210 0 90 $X=35690 $Y=2130
X355 64 M2_M1_CDNS_11 $T=37240 38080 0 0 $X=37160 $Y=37950
X356 73 M2_M1_CDNS_11 $T=41060 27730 0 0 $X=40980 $Y=27600
X357 63 M2_M1_CDNS_11 $T=43080 53380 0 0 $X=43000 $Y=53250
X358 7 M2_M1_CDNS_11 $T=47420 36740 0 0 $X=47340 $Y=36610
X359 49 M2_M1_CDNS_11 $T=47770 37090 0 0 $X=47690 $Y=36960
X360 67 M2_M1_CDNS_11 $T=50960 49840 0 90 $X=50830 $Y=49760
X361 47 M2_M1_CDNS_11 $T=51290 41540 0 90 $X=51160 $Y=41460
X362 65 M2_M1_CDNS_11 $T=51280 20630 0 0 $X=51200 $Y=20500
X363 70 M2_M1_CDNS_11 $T=51290 35200 0 0 $X=51210 $Y=35070
X364 60 M2_M1_CDNS_11 $T=51300 27960 0 0 $X=51220 $Y=27830
X365 72 M2_M1_CDNS_11 $T=51300 57100 0 0 $X=51220 $Y=56970
X366 57 M2_M1_CDNS_11 $T=59660 8330 0 0 $X=59580 $Y=8200
X367 71 M2_M1_CDNS_11 $T=59660 15640 0 0 $X=59580 $Y=15510
X368 69 M2_M1_CDNS_11 $T=59660 22940 0 0 $X=59580 $Y=22810
X369 54 M2_M1_CDNS_11 $T=59660 30310 0 0 $X=59580 $Y=30180
X370 49 M2_M1_CDNS_11 $T=59660 37620 0 0 $X=59580 $Y=37490
X371 55 M2_M1_CDNS_11 $T=59660 44940 0 0 $X=59580 $Y=44810
X372 53 M2_M1_CDNS_11 $T=59660 52270 0 0 $X=59580 $Y=52140
X373 67 M4_M3_CDNS_12 $T=32380 35710 0 90 $X=32130 $Y=35630
X374 68 M4_M3_CDNS_12 $T=33360 32510 0 90 $X=33110 $Y=32430
X375 55 M4_M3_CDNS_12 $T=33880 28620 0 0 $X=33800 $Y=28370
X376 53 M4_M3_CDNS_12 $T=34010 30140 0 0 $X=33930 $Y=29890
X377 54 M4_M3_CDNS_12 $T=34370 21060 0 0 $X=34290 $Y=20810
X378 69 M4_M3_CDNS_12 $T=36160 20250 0 0 $X=36080 $Y=20000
X379 71 M4_M3_CDNS_12 $T=36500 13950 0 0 $X=36420 $Y=13700
X380 72 M4_M3_CDNS_12 $T=37400 32460 0 0 $X=37320 $Y=32210
X381 65 M4_M3_CDNS_12 $T=37820 20120 0 0 $X=37740 $Y=19870
X382 71 M4_M3_CDNS_12 $T=40460 17040 0 90 $X=40210 $Y=16960
X383 65 M4_M3_CDNS_12 $T=40660 20120 0 90 $X=40410 $Y=20040
X384 57 M4_M3_CDNS_12 $T=40730 9730 0 90 $X=40480 $Y=9650
X385 60 M4_M3_CDNS_12 $T=40560 26320 0 0 $X=40480 $Y=26070
X386 72 M4_M3_CDNS_12 $T=42630 35130 0 90 $X=42380 $Y=35050
X387 7 M4_M3_CDNS_12 $T=47890 45870 0 0 $X=47810 $Y=45620
X388 6 M1_PO_CDNS_13 $T=1860 60810 0 0 $X=1760 $Y=60560
X389 6 M1_PO_CDNS_13 $T=1870 68120 0 0 $X=1770 $Y=67870
X390 4 M1_PO_CDNS_13 $T=2350 44590 0 90 $X=2100 $Y=44490
X391 3 M1_PO_CDNS_13 $T=3900 48300 0 90 $X=3650 $Y=48200
X392 2 M1_PO_CDNS_13 $T=3940 58210 0 90 $X=3690 $Y=58110
X393 10 M1_PO_CDNS_13 $T=6840 58120 0 90 $X=6590 $Y=58020
X394 6 M1_PO_CDNS_13 $T=12100 60800 0 0 $X=12000 $Y=60550
X395 6 M1_PO_CDNS_13 $T=12100 68120 0 0 $X=12000 $Y=67870
X396 6 M1_PO_CDNS_13 $T=22340 68120 0 0 $X=22240 $Y=67870
X397 6 M1_PO_CDNS_13 $T=22350 60800 0 0 $X=22250 $Y=60550
X398 6 M1_PO_CDNS_13 $T=32580 60800 0 0 $X=32480 $Y=60550
X399 6 M1_PO_CDNS_13 $T=32580 68120 0 0 $X=32480 $Y=67870
X400 52 M1_PO_CDNS_13 $T=33670 6150 0 90 $X=33420 $Y=6050
X401 6 M1_PO_CDNS_13 $T=40360 10220 0 90 $X=40110 $Y=10120
X402 6 M1_PO_CDNS_13 $T=40340 24940 0 0 $X=40240 $Y=24690
X403 6 M1_PO_CDNS_13 $T=40370 17590 0 0 $X=40270 $Y=17340
X404 7 M1_PO_CDNS_13 $T=46890 13630 0 0 $X=46790 $Y=13380
X405 7 M1_PO_CDNS_13 $T=46900 20740 0 0 $X=46800 $Y=20490
X406 7 M1_PO_CDNS_13 $T=46910 28080 0 0 $X=46810 $Y=27830
X407 6 M1_PO_CDNS_13 $T=47620 54480 0 90 $X=47370 $Y=54380
X408 6 M1_PO_CDNS_13 $T=47800 38230 0 90 $X=47550 $Y=38130
X409 6 M1_PO_CDNS_13 $T=47870 10240 0 0 $X=47770 $Y=9990
X410 6 M1_PO_CDNS_13 $T=47980 9490 0 0 $X=47880 $Y=9240
X411 6 M1_PO_CDNS_13 $T=48260 51950 0 90 $X=48010 $Y=51850
X412 6 M1_PO_CDNS_13 $T=48260 45130 0 0 $X=48160 $Y=44880
X413 6 M1_PO_CDNS_13 $T=48690 16910 0 0 $X=48590 $Y=16660
X414 6 M1_PO_CDNS_13 $T=48860 24230 0 0 $X=48760 $Y=23980
X415 6 M1_PO_CDNS_13 $T=48880 2280 0 0 $X=48780 $Y=2030
X416 56 M3_M2_CDNS_14 $T=14040 560 0 0 $X=13960 $Y=430
X417 59 M3_M2_CDNS_14 $T=22250 3160 0 0 $X=22170 $Y=3030
X418 56 M3_M2_CDNS_14 $T=23920 6540 0 0 $X=23840 $Y=6410
X419 48 M3_M2_CDNS_14 $T=25520 48970 0 0 $X=25440 $Y=48840
X420 64 M3_M2_CDNS_14 $T=27740 16660 0 0 $X=27660 $Y=16530
X421 51 M3_M2_CDNS_14 $T=28010 24010 0 0 $X=27930 $Y=23880
X422 72 M3_M2_CDNS_14 $T=31460 30680 0 90 $X=31330 $Y=30600
X423 48 M3_M2_CDNS_14 $T=32190 54030 0 0 $X=32110 $Y=53900
X424 68 M3_M2_CDNS_14 $T=36910 32510 0 0 $X=36830 $Y=32380
X425 68 M3_M2_CDNS_14 $T=37470 13030 0 0 $X=37390 $Y=12900
X426 73 M3_M2_CDNS_14 $T=37590 8380 0 90 $X=37460 $Y=8300
X427 73 M3_M2_CDNS_14 $T=38080 28430 0 0 $X=38000 $Y=28300
X428 49 M3_M2_CDNS_14 $T=39590 33870 0 0 $X=39510 $Y=33740
X429 67 M3_M2_CDNS_14 $T=40110 35670 0 90 $X=39980 $Y=35590
X430 70 M3_M2_CDNS_14 $T=42020 34330 0 0 $X=41940 $Y=34200
X431 55 M3_M2_CDNS_14 $T=45640 37660 0 0 $X=45560 $Y=37530
X432 6 M3_M2_CDNS_14 $T=47780 30450 0 0 $X=47700 $Y=30320
X433 6 M3_M2_CDNS_14 $T=47810 35930 0 0 $X=47730 $Y=35800
X434 65 M3_M2_CDNS_14 $T=48170 20860 0 0 $X=48090 $Y=20730
X435 60 M3_M2_CDNS_14 $T=48180 28260 0 0 $X=48100 $Y=28130
X436 7 M3_M2_CDNS_14 $T=48350 54060 0 0 $X=48270 $Y=53930
X437 71 M3_M2_CDNS_14 $T=48430 15830 0 0 $X=48350 $Y=15700
X438 72 M3_M2_CDNS_14 $T=49580 57720 0 90 $X=49450 $Y=57640
X439 57 M3_M2_CDNS_14 $T=50600 8490 0 0 $X=50520 $Y=8360
X440 6 M1_PO_CDNS_15 $T=47780 31470 0 0 $X=47680 $Y=31220
X441 7 M1_PO_CDNS_16 $T=47950 48930 0 0 $X=47850 $Y=48810
X442 6 M2_M1_CDNS_17 $T=47780 31470 0 0 $X=47700 $Y=31220
X443 1 5 2 3 4 9 14 13 10 50
+ 15 46 62 48 68 64 51 63 251 260
+ 231 228 214 224 218 288 249 250 253 313
+ 314 307 275 232 279 290 266 317 318 278
+ 216 289 277 293 296 219 300 262 316 261 multiplier $T=1090 33260 0 0 $X=750 $Y=33040
X444 56 19 9 5 8 64 48 52 57 71
+ 54 49 55 53 63 51 62 69 68 50
+ 46 59 58 18 72 70 47 67 73 61
+ 65 60 66 74 95 112 111 110 109 115
+ 114 121 120 119 118 103 102 105 104 141
+ 211 107 106 97 96 99 98 101 100 108
+ 113 130 139 140 158 159 176 185 190 191
+ 194 212 213 760 761 762 763 10badder $T=-50390 53780 1 0 $X=-110 $Y=0
X445 9 7 5 6 1 11 90 86 91 87
+ 506 88 508 84 85 89 92 ph1p3_MSDFF $T=1140 62320 0 0 $X=1140 $Y=58560
X446 9 7 5 6 2 12 81 77 82 78
+ 503 79 505 75 76 80 83 ph1p3_MSDFF $T=1140 69640 0 0 $X=1140 $Y=65880
X447 9 7 5 6 14 17 345 341 346 342
+ 692 343 694 339 340 344 347 ph1p3_MSDFF $T=11380 62320 0 0 $X=11380 $Y=58560
X448 9 7 5 6 10 16 336 332 337 333
+ 689 334 691 330 331 335 338 ph1p3_MSDFF $T=11380 69640 0 0 $X=11380 $Y=65880
X449 9 7 5 6 13 21 363 359 364 360
+ 698 361 700 357 358 362 365 ph1p3_MSDFF $T=21620 62320 0 0 $X=21620 $Y=58560
X450 9 7 5 6 3 20 354 350 355 351
+ 695 352 697 348 349 353 356 ph1p3_MSDFF $T=21620 69640 0 0 $X=21620 $Y=65880
X451 9 7 5 6 15 22 381 377 382 378
+ 704 379 706 375 376 380 383 ph1p3_MSDFF $T=31860 62320 0 0 $X=31860 $Y=58560
X452 9 7 5 6 4 23 372 368 373 369
+ 701 370 703 366 367 371 374 ph1p3_MSDFF $T=31860 69640 0 0 $X=31860 $Y=65880
X453 9 7 5 6 66 58 408 404 409 405
+ 713 406 715 402 403 407 410 ph1p3_MSDFF $T=37920 11080 0 0 $X=37920 $Y=7320
X454 9 7 5 6 59 56 399 395 400 396
+ 710 397 712 393 394 398 401 ph1p3_MSDFF $T=37920 18400 0 0 $X=37920 $Y=14640
X455 9 7 5 6 73 52 390 386 391 387
+ 707 388 709 384 385 389 392 ph1p3_MSDFF $T=37920 25720 0 0 $X=37920 $Y=21960
X456 9 7 5 6 24 25 480 476 481 477
+ 737 478 739 474 475 479 482 ph1p3_MSDFF $T=48160 3760 0 0 $X=48160 $Y=0
X457 9 7 5 6 61 57 471 467 472 468
+ 734 469 736 465 466 470 473 ph1p3_MSDFF $T=48160 11080 0 0 $X=48160 $Y=7320
X458 9 7 5 6 65 71 462 458 463 459
+ 731 460 733 456 457 461 464 ph1p3_MSDFF $T=48160 18400 0 0 $X=48160 $Y=14640
X459 9 7 5 6 60 69 453 449 454 450
+ 728 451 730 447 448 452 455 ph1p3_MSDFF $T=48160 25720 0 0 $X=48160 $Y=21960
X460 9 7 5 6 70 54 444 440 445 441
+ 725 442 727 438 439 443 446 ph1p3_MSDFF $T=48160 33040 0 0 $X=48160 $Y=29280
X461 9 7 5 6 47 49 435 431 436 432
+ 722 433 724 429 430 434 437 ph1p3_MSDFF $T=48160 40360 0 0 $X=48160 $Y=36600
X462 9 7 5 6 67 55 426 422 427 423
+ 719 424 721 420 421 425 428 ph1p3_MSDFF $T=48160 47680 0 0 $X=48160 $Y=43920
X463 9 7 5 6 72 53 417 413 418 414
+ 716 415 718 411 412 416 419 ph1p3_MSDFF $T=48160 55000 0 0 $X=48160 $Y=51240
X464 9 5 cellTmpl_CDNS_49 $T=47620 54900 1 0 $X=47500 $Y=51240
X465 25 57 9 5 36 34 501 502 758 759
+ 788 789 MUX_2to1___2X_ph2p2 $T=58160 11120 1 0 $X=58160 $Y=7320
X466 25 58 9 5 37 29 499 500 756 757
+ 786 787 MUX_2to1___2X_ph2p2 $T=58160 11080 0 0 $X=58160 $Y=11080
X467 25 71 9 5 38 26 497 498 754 755
+ 784 785 MUX_2to1___2X_ph2p2 $T=58160 18440 1 0 $X=58160 $Y=14640
X468 25 56 9 5 39 31 495 496 752 753
+ 782 783 MUX_2to1___2X_ph2p2 $T=58160 18400 0 0 $X=58160 $Y=18400
X469 25 69 9 5 40 32 493 494 750 751
+ 780 781 MUX_2to1___2X_ph2p2 $T=58160 25760 1 0 $X=58160 $Y=21960
X470 25 52 9 5 41 35 491 492 748 749
+ 778 779 MUX_2to1___2X_ph2p2 $T=58160 25720 0 0 $X=58160 $Y=25720
X471 25 54 9 5 42 28 489 490 746 747
+ 776 777 MUX_2to1___2X_ph2p2 $T=58160 33080 1 0 $X=58160 $Y=29280
X472 25 49 9 5 43 33 487 488 744 745
+ 774 775 MUX_2to1___2X_ph2p2 $T=58160 40400 1 0 $X=58160 $Y=36600
X473 25 55 9 5 44 30 485 486 742 743
+ 772 773 MUX_2to1___2X_ph2p2 $T=58160 47720 1 0 $X=58160 $Y=43920
X474 25 53 9 5 45 27 483 484 740 741
+ 770 771 MUX_2to1___2X_ph2p2 $T=58160 55040 1 0 $X=58160 $Y=51240
M0 87 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=59450 $dt=1
M1 90 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=64750 $dt=1
M2 78 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=66770 $dt=1
M3 84 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3250 $Y=64780 $dt=1
M4 85 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=59420 $dt=1
M5 76 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=66740 $dt=1
M6 86 7 1 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4430 $Y=64780 $dt=1
M7 91 7 506 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=59660 $dt=1
M8 82 7 503 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=66980 $dt=1
M9 88 86 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5630 $Y=64690 $dt=1
M10 506 11 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=59450 $dt=1
M11 503 12 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=66770 $dt=1
M12 88 87 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6870 $Y=64700 $dt=1
M13 89 90 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=59420 $dt=1
M14 80 81 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=66740 $dt=1
M15 508 88 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8120 $Y=64750 $dt=1
M16 91 90 88 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=59660 $dt=1
M17 82 81 79 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=66980 $dt=1
M18 92 90 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9450 $Y=64780 $dt=1
M19 11 91 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=59450 $dt=1
M20 12 82 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=66770 $dt=1
M21 86 90 508 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=10630 $Y=64780 $dt=1
M22 342 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=59450 $dt=1
M23 345 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=64750 $dt=1
M24 333 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=66770 $dt=1
M25 339 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13490 $Y=64780 $dt=1
M26 340 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=59420 $dt=1
M27 331 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=66740 $dt=1
M28 341 7 14 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=14670 $Y=64780 $dt=1
M29 346 7 692 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=59660 $dt=1
M30 337 7 689 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=66980 $dt=1
M31 343 341 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=15870 $Y=64690 $dt=1
M32 692 17 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=59450 $dt=1
M33 689 16 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=66770 $dt=1
M34 343 342 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17110 $Y=64700 $dt=1
M35 344 345 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=59420 $dt=1
M36 335 336 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=66740 $dt=1
M37 694 343 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18360 $Y=64750 $dt=1
M38 346 345 343 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=59660 $dt=1
M39 337 336 334 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=66980 $dt=1
M40 347 345 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=19690 $Y=64780 $dt=1
M41 17 346 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=59450 $dt=1
M42 16 337 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=66770 $dt=1
M43 341 345 694 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=20870 $Y=64780 $dt=1
M44 360 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=59450 $dt=1
M45 363 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=64750 $dt=1
M46 351 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=66770 $dt=1
M47 357 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=23730 $Y=64780 $dt=1
M48 358 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=59420 $dt=1
M49 349 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=66740 $dt=1
M50 359 7 13 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=24910 $Y=64780 $dt=1
M51 364 7 698 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=59660 $dt=1
M52 355 7 695 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=66980 $dt=1
M53 361 359 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26110 $Y=64690 $dt=1
M54 698 21 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=59450 $dt=1
M55 695 20 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=66770 $dt=1
M56 361 360 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27350 $Y=64700 $dt=1
M57 362 363 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=59420 $dt=1
M58 353 354 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=66740 $dt=1
M59 700 361 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28600 $Y=64750 $dt=1
M60 364 363 361 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=59660 $dt=1
M61 355 354 352 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=66980 $dt=1
M62 365 363 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=29930 $Y=64780 $dt=1
M63 21 364 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=59450 $dt=1
M64 20 355 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=66770 $dt=1
M65 359 363 700 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31110 $Y=64780 $dt=1
M66 378 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=59450 $dt=1
M67 381 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=64750 $dt=1
M68 369 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=66770 $dt=1
M69 375 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=33970 $Y=64780 $dt=1
M70 376 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=59420 $dt=1
M71 367 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=66740 $dt=1
M72 377 7 15 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35150 $Y=64780 $dt=1
M73 382 7 704 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=59660 $dt=1
M74 373 7 701 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=66980 $dt=1
M75 379 377 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36350 $Y=64690 $dt=1
M76 704 22 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=37440 $Y=59450 $dt=1
M77 701 23 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=37440 $Y=66770 $dt=1
M78 379 378 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37590 $Y=64700 $dt=1
M79 405 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=8210 $dt=1
M80 408 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=13510 $dt=1
M81 396 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=15530 $dt=1
M82 399 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=20830 $dt=1
M83 387 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=22850 $dt=1
M84 390 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=28150 $dt=1
M85 380 381 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=38770 $Y=59420 $dt=1
M86 371 372 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=38770 $Y=66740 $dt=1
M87 706 379 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=38840 $Y=64750 $dt=1
M88 382 381 379 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=39950 $Y=59660 $dt=1
M89 373 372 370 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=39950 $Y=66980 $dt=1
M90 402 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=13540 $dt=1
M91 393 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=20860 $dt=1
M92 384 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=40030 $Y=28180 $dt=1
M93 383 381 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40170 $Y=64780 $dt=1
M94 403 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=41030 $Y=8180 $dt=1
M95 394 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=15500 $dt=1
M96 385 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=22820 $dt=1
M97 404 7 66 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=13540 $dt=1
M98 395 7 59 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=20860 $dt=1
M99 386 7 73 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=41210 $Y=28180 $dt=1
M100 22 382 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=41240 $Y=59450 $dt=1
M101 23 373 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=41240 $Y=66770 $dt=1
M102 377 381 706 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41350 $Y=64780 $dt=1
M103 409 7 713 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=42210 $Y=8420 $dt=1
M104 400 7 710 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=15740 $dt=1
M105 391 7 707 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=23060 $dt=1
M106 406 404 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=13450 $dt=1
M107 397 395 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=20770 $dt=1
M108 388 386 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42410 $Y=28090 $dt=1
M109 713 58 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=43500 $Y=8210 $dt=1
M110 710 56 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=15530 $dt=1
M111 707 52 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=22850 $dt=1
M112 406 405 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=13460 $dt=1
M113 397 396 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=20780 $dt=1
M114 388 387 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43650 $Y=28100 $dt=1
M115 407 408 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=44830 $Y=8180 $dt=1
M116 398 399 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=15500 $dt=1
M117 389 390 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=22820 $dt=1
M118 715 406 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=13510 $dt=1
M119 712 397 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=20830 $dt=1
M120 709 388 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=44900 $Y=28150 $dt=1
M121 409 408 406 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=46010 $Y=8420 $dt=1
M122 400 399 397 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=15740 $dt=1
M123 391 390 388 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=23060 $dt=1
M124 410 408 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=13540 $dt=1
M125 401 399 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=20860 $dt=1
M126 392 390 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=46230 $Y=28180 $dt=1
M127 58 409 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=47300 $Y=8210 $dt=1
M128 56 400 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=15530 $dt=1
M129 52 391 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=22850 $dt=1
M130 404 408 715 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=13540 $dt=1
M131 395 399 712 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=20860 $dt=1
M132 386 390 709 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=47410 $Y=28180 $dt=1
M133 477 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=890 $dt=1
M134 480 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=6190 $dt=1
M135 468 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=8210 $dt=1
M136 471 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=13510 $dt=1
M137 459 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=15530 $dt=1
M138 462 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=20830 $dt=1
M139 450 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=22850 $dt=1
M140 453 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=28150 $dt=1
M141 441 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=30170 $dt=1
M142 444 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=35470 $dt=1
M143 432 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=37490 $dt=1
M144 435 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=42790 $dt=1
M145 423 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=44810 $dt=1
M146 426 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=50110 $dt=1
M147 414 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=52130 $dt=1
M148 417 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=57430 $dt=1
M149 474 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=6220 $dt=1
M150 465 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=13540 $dt=1
M151 456 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=20860 $dt=1
M152 447 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=28180 $dt=1
M153 438 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=35500 $dt=1
M154 429 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=42820 $dt=1
M155 420 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=50140 $dt=1
M156 411 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=50270 $Y=57460 $dt=1
M157 475 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=51270 $Y=860 $dt=1
M158 466 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=8180 $dt=1
M159 457 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=15500 $dt=1
M160 448 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=22820 $dt=1
M161 439 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=30140 $dt=1
M162 430 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=37460 $dt=1
M163 421 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=44780 $dt=1
M164 412 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=52100 $dt=1
M165 476 7 24 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=6220 $dt=1
M166 467 7 61 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=13540 $dt=1
M167 458 7 65 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=20860 $dt=1
M168 449 7 60 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=28180 $dt=1
M169 440 7 70 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=35500 $dt=1
M170 431 7 47 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=42820 $dt=1
M171 422 7 67 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=50140 $dt=1
M172 413 7 72 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=51450 $Y=57460 $dt=1
M173 481 7 737 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=52450 $Y=1100 $dt=1
M174 472 7 734 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=8420 $dt=1
M175 463 7 731 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=15740 $dt=1
M176 454 7 728 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=23060 $dt=1
M177 445 7 725 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=30380 $dt=1
M178 436 7 722 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=37700 $dt=1
M179 427 7 719 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=45020 $dt=1
M180 418 7 716 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=52340 $dt=1
M181 478 476 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=6130 $dt=1
M182 469 467 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=13450 $dt=1
M183 460 458 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=20770 $dt=1
M184 451 449 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=28090 $dt=1
M185 442 440 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=35410 $dt=1
M186 433 431 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=42730 $dt=1
M187 424 422 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=50050 $dt=1
M188 415 413 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=52650 $Y=57370 $dt=1
M189 737 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=53740 $Y=890 $dt=1
M190 734 57 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=8210 $dt=1
M191 731 71 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=15530 $dt=1
M192 728 69 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=22850 $dt=1
M193 725 54 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=30170 $dt=1
M194 722 49 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=37490 $dt=1
M195 719 55 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=44810 $dt=1
M196 716 53 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=52130 $dt=1
M197 478 477 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=6140 $dt=1
M198 469 468 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=13460 $dt=1
M199 460 459 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=20780 $dt=1
M200 451 450 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=28100 $dt=1
M201 442 441 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=35420 $dt=1
M202 433 432 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=42740 $dt=1
M203 424 423 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=50060 $dt=1
M204 415 414 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=53890 $Y=57380 $dt=1
M205 479 480 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=55070 $Y=860 $dt=1
M206 470 471 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=8180 $dt=1
M207 461 462 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=15500 $dt=1
M208 452 453 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=22820 $dt=1
M209 443 444 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=30140 $dt=1
M210 434 435 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=37460 $dt=1
M211 425 426 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=44780 $dt=1
M212 416 417 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=52100 $dt=1
M213 739 478 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=6190 $dt=1
M214 736 469 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=13510 $dt=1
M215 733 460 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=20830 $dt=1
M216 730 451 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=28150 $dt=1
M217 727 442 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=35470 $dt=1
M218 724 433 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=42790 $dt=1
M219 721 424 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=50110 $dt=1
M220 718 415 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=55140 $Y=57430 $dt=1
M221 481 480 478 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=56250 $Y=1100 $dt=1
M222 472 471 469 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=8420 $dt=1
M223 463 462 460 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=15740 $dt=1
M224 454 453 451 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=23060 $dt=1
M225 445 444 442 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=30380 $dt=1
M226 436 435 433 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=37700 $dt=1
M227 427 426 424 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=45020 $dt=1
M228 418 417 415 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=52340 $dt=1
M229 482 480 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=6220 $dt=1
M230 473 471 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=13540 $dt=1
M231 464 462 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=20860 $dt=1
M232 455 453 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=28180 $dt=1
M233 446 444 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=35500 $dt=1
M234 437 435 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=42820 $dt=1
M235 428 426 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=50140 $dt=1
M236 419 417 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=56470 $Y=57460 $dt=1
M237 25 481 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=57540 $Y=890 $dt=1
M238 57 472 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=8210 $dt=1
M239 71 463 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=15530 $dt=1
M240 69 454 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=22850 $dt=1
M241 54 445 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=30170 $dt=1
M242 49 436 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=37490 $dt=1
M243 55 427 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=44810 $dt=1
M244 53 418 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=52130 $dt=1
M245 476 480 739 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=6220 $dt=1
M246 467 471 736 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=13540 $dt=1
M247 458 462 733 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=20860 $dt=1
M248 449 453 730 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=28180 $dt=1
M249 440 444 727 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=35500 $dt=1
M250 431 435 724 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=42820 $dt=1
M251 422 426 721 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=50140 $dt=1
M252 413 417 718 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=57650 $Y=57460 $dt=1
M253 501 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=8270 $dt=1
M254 499 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=13450 $dt=1
M255 497 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=15590 $dt=1
M256 495 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=20770 $dt=1
M257 493 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=22910 $dt=1
M258 491 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=28090 $dt=1
M259 489 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=30230 $dt=1
M260 487 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=37550 $dt=1
M261 485 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=44870 $dt=1
M262 483 25 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=52190 $dt=1
M263 788 57 502 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=8060 $dt=1
M264 786 58 500 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=13180 $dt=1
M265 784 71 498 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=15380 $dt=1
M266 782 56 496 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=20500 $dt=1
M267 780 69 494 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=22700 $dt=1
M268 778 52 492 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=27820 $dt=1
M269 776 54 490 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=30020 $dt=1
M270 774 49 488 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=37340 $dt=1
M271 772 55 486 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=44660 $dt=1
M272 770 53 484 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=51980 $dt=1
M273 9 25 788 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=8060 $dt=1
M274 9 25 786 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=13180 $dt=1
M275 9 25 784 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=15380 $dt=1
M276 9 25 782 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=20500 $dt=1
M277 9 25 780 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=22700 $dt=1
M278 9 25 778 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=27820 $dt=1
M279 9 25 776 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=30020 $dt=1
M280 9 25 774 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=37340 $dt=1
M281 9 25 772 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=44660 $dt=1
M282 9 25 770 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=51980 $dt=1
M283 789 501 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=8130 $dt=1
M284 787 499 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=13110 $dt=1
M285 785 497 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=15450 $dt=1
M286 783 495 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=20430 $dt=1
M287 781 493 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=22770 $dt=1
M288 779 491 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=27750 $dt=1
M289 777 489 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=30090 $dt=1
M290 775 487 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=37410 $dt=1
M291 773 485 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=44730 $dt=1
M292 771 483 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=52050 $dt=1
M293 502 36 789 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=8130 $dt=1
M294 500 37 787 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=13110 $dt=1
M295 498 38 785 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=15450 $dt=1
M296 496 39 783 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=20430 $dt=1
M297 494 40 781 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=22770 $dt=1
M298 492 41 779 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=27750 $dt=1
M299 490 42 777 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=30090 $dt=1
M300 488 43 775 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=37410 $dt=1
M301 486 44 773 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=44730 $dt=1
M302 484 45 771 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=52050 $dt=1
M303 34 502 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=8120 $dt=1
M304 29 500 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=13120 $dt=1
M305 26 498 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=15440 $dt=1
M306 31 496 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=20440 $dt=1
M307 32 494 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=22760 $dt=1
M308 35 492 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=27760 $dt=1
M309 28 490 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=30080 $dt=1
M310 33 488 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=37400 $dt=1
M311 30 486 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=44720 $dt=1
M312 27 484 9 9 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=52040 $dt=1
.ends ph2p2_processing_element

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p3_Matrix_vector_Multiplication              *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p3_Matrix_vector_Multiplication 109 107 108 100 104 111 114 113 110 106
+ 92 90 91 87 88 94 97 96 93 89
+ 79 77 78 74 75 81 84 83 80 76
+ 53 51 52 44 47 56 60 59 55 49
+ 101 105 102 103 50 54 58 61 46 112
+ 95 82 57 1 115 116 98 99 85 86
+ 62 63 73 72 71 70 68 66 64 69
+ 67 65 118 121 124 119 123 117 125 126
+ 122 120 45 48
** N=2230 EP=84 FDC=6648
X0 1 M3_M2_CDNS_1 $T=47980 58060 0 90 $X=47730 $Y=57980
X1 1 M3_M2_CDNS_1 $T=47980 131280 0 90 $X=47730 $Y=131200
X2 1 M3_M2_CDNS_1 $T=47980 204490 0 90 $X=47730 $Y=204410
X3 2 M3_M2_CDNS_1 $T=63820 31300 0 0 $X=63740 $Y=31050
X4 2 M3_M2_CDNS_1 $T=63820 71930 0 0 $X=63740 $Y=71680
X5 3 M3_M2_CDNS_1 $T=63820 104520 0 0 $X=63740 $Y=104270
X6 3 M3_M2_CDNS_1 $T=63820 145150 0 0 $X=63740 $Y=144900
X7 4 M3_M2_CDNS_1 $T=63820 177730 0 0 $X=63740 $Y=177480
X8 4 M3_M2_CDNS_1 $T=63820 218360 0 0 $X=63740 $Y=218110
X9 5 M3_M2_CDNS_1 $T=63850 23980 0 0 $X=63770 $Y=23730
X10 6 M3_M2_CDNS_1 $T=63850 97200 0 0 $X=63770 $Y=96950
X11 7 M3_M2_CDNS_1 $T=63850 170410 0 0 $X=63770 $Y=170160
X12 8 M3_M2_CDNS_1 $T=63890 27300 0 0 $X=63810 $Y=27050
X13 9 M3_M2_CDNS_1 $T=63890 100520 0 0 $X=63810 $Y=100270
X14 10 M3_M2_CDNS_1 $T=63890 173730 0 0 $X=63810 $Y=173480
X15 1 M2_M1_CDNS_2 $T=47980 58060 0 90 $X=47730 $Y=57980
X16 1 M2_M1_CDNS_2 $T=47980 131280 0 90 $X=47730 $Y=131200
X17 1 M2_M1_CDNS_2 $T=47980 204490 0 90 $X=47730 $Y=204410
X18 2 M2_M1_CDNS_2 $T=63820 31300 0 0 $X=63740 $Y=31050
X19 2 M2_M1_CDNS_2 $T=63820 71930 0 0 $X=63740 $Y=71680
X20 3 M2_M1_CDNS_2 $T=63820 104520 0 0 $X=63740 $Y=104270
X21 3 M2_M1_CDNS_2 $T=63820 145150 0 0 $X=63740 $Y=144900
X22 4 M2_M1_CDNS_2 $T=63820 177730 0 0 $X=63740 $Y=177480
X23 4 M2_M1_CDNS_2 $T=63820 218360 0 0 $X=63740 $Y=218110
X24 5 M2_M1_CDNS_2 $T=63850 23980 0 0 $X=63770 $Y=23730
X25 6 M2_M1_CDNS_2 $T=63850 97200 0 0 $X=63770 $Y=96950
X26 7 M2_M1_CDNS_2 $T=63850 170410 0 0 $X=63770 $Y=170160
X27 8 M2_M1_CDNS_2 $T=63890 27300 0 0 $X=63810 $Y=27050
X28 9 M2_M1_CDNS_2 $T=63890 100520 0 0 $X=63810 $Y=100270
X29 10 M2_M1_CDNS_2 $T=63890 173730 0 0 $X=63810 $Y=173480
X30 11 M5_M4_CDNS_3 $T=9410 93400 0 0 $X=9330 $Y=93270
X31 12 M5_M4_CDNS_3 $T=9410 166620 0 0 $X=9330 $Y=166490
X32 13 M5_M4_CDNS_3 $T=9410 239830 0 0 $X=9330 $Y=239700
X33 14 M5_M4_CDNS_3 $T=9820 94000 0 0 $X=9740 $Y=93870
X34 15 M5_M4_CDNS_3 $T=9820 167220 0 0 $X=9740 $Y=167090
X35 16 M5_M4_CDNS_3 $T=9820 240430 0 0 $X=9740 $Y=240300
X36 17 M5_M4_CDNS_3 $T=25120 73790 0 0 $X=25040 $Y=73660
X37 18 M5_M4_CDNS_3 $T=25120 147010 0 0 $X=25040 $Y=146880
X38 19 M5_M4_CDNS_3 $T=25120 220220 0 0 $X=25040 $Y=220090
X39 20 M5_M4_CDNS_3 $T=28450 130040 0 0 $X=28370 $Y=129910
X40 21 M5_M4_CDNS_3 $T=28450 203260 0 0 $X=28370 $Y=203130
X41 22 M5_M4_CDNS_3 $T=28450 276470 0 0 $X=28370 $Y=276340
X42 17 M5_M4_CDNS_3 $T=30670 73840 0 0 $X=30590 $Y=73710
X43 18 M5_M4_CDNS_3 $T=30670 147060 0 0 $X=30590 $Y=146930
X44 19 M5_M4_CDNS_3 $T=30670 220270 0 0 $X=30590 $Y=220140
X45 17 M5_M4_CDNS_3 $T=35390 130710 0 0 $X=35310 $Y=130580
X46 18 M5_M4_CDNS_3 $T=35390 203930 0 0 $X=35310 $Y=203800
X47 19 M5_M4_CDNS_3 $T=35390 277140 0 0 $X=35310 $Y=277010
X48 23 M5_M4_CDNS_3 $T=55470 70970 0 90 $X=55340 $Y=70890
X49 24 M5_M4_CDNS_3 $T=55470 144190 0 90 $X=55340 $Y=144110
X50 25 M5_M4_CDNS_3 $T=55470 217400 0 90 $X=55340 $Y=217320
X51 8 M5_M4_CDNS_3 $T=56490 100610 0 90 $X=56360 $Y=100530
X52 9 M5_M4_CDNS_3 $T=56490 173830 0 90 $X=56360 $Y=173750
X53 10 M5_M4_CDNS_3 $T=56490 247040 0 90 $X=56360 $Y=246960
X54 5 M5_M4_CDNS_3 $T=56560 97140 0 0 $X=56480 $Y=97010
X55 6 M5_M4_CDNS_3 $T=56560 170360 0 0 $X=56480 $Y=170230
X56 7 M5_M4_CDNS_3 $T=56560 243570 0 0 $X=56480 $Y=243440
X57 26 M5_M4_CDNS_3 $T=57090 92750 0 0 $X=57010 $Y=92620
X58 27 M5_M4_CDNS_3 $T=57090 165970 0 0 $X=57010 $Y=165840
X59 28 M5_M4_CDNS_3 $T=57090 239180 0 0 $X=57010 $Y=239050
X60 29 M5_M4_CDNS_3 $T=57150 110830 0 0 $X=57070 $Y=110700
X61 30 M5_M4_CDNS_3 $T=57150 184050 0 0 $X=57070 $Y=183920
X62 31 M5_M4_CDNS_3 $T=57150 257260 0 0 $X=57070 $Y=257130
X63 32 M5_M4_CDNS_3 $T=57170 125430 0 0 $X=57090 $Y=125300
X64 33 M5_M4_CDNS_3 $T=57170 198650 0 0 $X=57090 $Y=198520
X65 34 M5_M4_CDNS_3 $T=57170 271860 0 0 $X=57090 $Y=271730
X66 35 M5_M4_CDNS_3 $T=57200 118260 0 0 $X=57120 $Y=118130
X67 36 M5_M4_CDNS_3 $T=57200 191480 0 0 $X=57120 $Y=191350
X68 37 M5_M4_CDNS_3 $T=57200 264690 0 0 $X=57120 $Y=264560
X69 2 M5_M4_CDNS_3 $T=57550 103260 0 0 $X=57470 $Y=103130
X70 3 M5_M4_CDNS_3 $T=57550 176480 0 0 $X=57470 $Y=176350
X71 4 M5_M4_CDNS_3 $T=57550 249690 0 0 $X=57470 $Y=249560
X72 4 M5_M4_CDNS_3 $T=62210 216190 0 90 $X=62080 $Y=216110
X73 3 M5_M4_CDNS_3 $T=62240 142980 0 90 $X=62110 $Y=142900
X74 2 M5_M4_CDNS_3 $T=62300 69760 0 90 $X=62170 $Y=69680
X75 32 M5_M4_CDNS_3 $T=62650 125410 0 0 $X=62570 $Y=125280
X76 33 M5_M4_CDNS_3 $T=62650 198630 0 0 $X=62570 $Y=198500
X77 34 M5_M4_CDNS_3 $T=62740 271840 0 0 $X=62660 $Y=271710
X78 29 M5_M4_CDNS_3 $T=62750 111060 0 0 $X=62670 $Y=110930
X79 30 M5_M4_CDNS_3 $T=62750 184280 0 0 $X=62670 $Y=184150
X80 31 M5_M4_CDNS_3 $T=62750 257490 0 0 $X=62670 $Y=257360
X81 35 M5_M4_CDNS_3 $T=62760 118220 0 0 $X=62680 $Y=118090
X82 36 M5_M4_CDNS_3 $T=62760 191440 0 0 $X=62680 $Y=191310
X83 37 M5_M4_CDNS_3 $T=62760 264650 0 0 $X=62680 $Y=264520
X84 11 M3_M2_CDNS_4 $T=11150 139470 0 90 $X=10900 $Y=139390
X85 12 M3_M2_CDNS_4 $T=11150 212690 0 90 $X=10900 $Y=212610
X86 13 M3_M2_CDNS_4 $T=11150 285900 0 90 $X=10900 $Y=285820
X87 14 M3_M2_CDNS_4 $T=16950 140010 0 180 $X=16870 $Y=139760
X88 15 M3_M2_CDNS_4 $T=16950 213230 0 180 $X=16870 $Y=212980
X89 16 M3_M2_CDNS_4 $T=16950 286440 0 180 $X=16870 $Y=286190
X90 20 M3_M2_CDNS_4 $T=31680 139470 0 90 $X=31430 $Y=139390
X91 21 M3_M2_CDNS_4 $T=31680 212690 0 90 $X=31430 $Y=212610
X92 22 M3_M2_CDNS_4 $T=31680 285900 0 90 $X=31430 $Y=285820
X93 17 M3_M2_CDNS_4 $T=41970 139470 0 90 $X=41720 $Y=139390
X94 18 M3_M2_CDNS_4 $T=41970 212690 0 90 $X=41720 $Y=212610
X95 19 M3_M2_CDNS_4 $T=41970 285900 0 90 $X=41720 $Y=285820
X96 29 M3_M2_CDNS_4 $T=51030 71710 0 0 $X=50950 $Y=71460
X97 30 M3_M2_CDNS_4 $T=51030 144930 0 0 $X=50950 $Y=144680
X98 31 M3_M2_CDNS_4 $T=51030 218140 0 0 $X=50950 $Y=217890
X99 35 M3_M2_CDNS_4 $T=51420 72540 0 0 $X=51340 $Y=72290
X100 36 M3_M2_CDNS_4 $T=51420 145760 0 0 $X=51340 $Y=145510
X101 37 M3_M2_CDNS_4 $T=51420 218970 0 0 $X=51340 $Y=218720
X102 32 M3_M2_CDNS_4 $T=54350 80260 0 0 $X=54270 $Y=80010
X103 33 M3_M2_CDNS_4 $T=54350 153480 0 0 $X=54270 $Y=153230
X104 34 M3_M2_CDNS_4 $T=54350 226690 0 0 $X=54270 $Y=226440
X105 4 M4_M3_CDNS_5 $T=62210 216190 0 90 $X=61960 $Y=216110
X106 3 M4_M3_CDNS_5 $T=62240 142980 0 90 $X=61990 $Y=142900
X107 2 M4_M3_CDNS_5 $T=62300 69760 0 90 $X=62050 $Y=69680
X108 32 M4_M3_CDNS_5 $T=62650 125410 0 0 $X=62570 $Y=125160
X109 33 M4_M3_CDNS_5 $T=62650 198630 0 0 $X=62570 $Y=198380
X110 2 M4_M3_CDNS_5 $T=62740 103290 0 0 $X=62660 $Y=103040
X111 3 M4_M3_CDNS_5 $T=62740 176510 0 0 $X=62660 $Y=176260
X112 4 M4_M3_CDNS_5 $T=62740 249720 0 0 $X=62660 $Y=249470
X113 34 M4_M3_CDNS_5 $T=62740 271840 0 0 $X=62660 $Y=271590
X114 38 M4_M3_CDNS_5 $T=62750 87190 0 0 $X=62670 $Y=86940
X115 29 M4_M3_CDNS_5 $T=62750 111060 0 0 $X=62670 $Y=110810
X116 39 M4_M3_CDNS_5 $T=62750 160410 0 0 $X=62670 $Y=160160
X117 30 M4_M3_CDNS_5 $T=62750 184280 0 0 $X=62670 $Y=184030
X118 40 M4_M3_CDNS_5 $T=62750 233620 0 0 $X=62670 $Y=233370
X119 31 M4_M3_CDNS_5 $T=62750 257490 0 0 $X=62670 $Y=257240
X120 41 M4_M3_CDNS_5 $T=62760 88540 0 0 $X=62680 $Y=88290
X121 26 M4_M3_CDNS_5 $T=62760 94470 0 0 $X=62680 $Y=94220
X122 5 M4_M3_CDNS_5 $T=62760 95900 0 0 $X=62680 $Y=95650
X123 8 M4_M3_CDNS_5 $T=62760 101860 0 0 $X=62680 $Y=101610
X124 35 M4_M3_CDNS_5 $T=62760 118220 0 0 $X=62680 $Y=117970
X125 42 M4_M3_CDNS_5 $T=62760 161760 0 0 $X=62680 $Y=161510
X126 27 M4_M3_CDNS_5 $T=62760 167690 0 0 $X=62680 $Y=167440
X127 6 M4_M3_CDNS_5 $T=62760 169120 0 0 $X=62680 $Y=168870
X128 9 M4_M3_CDNS_5 $T=62760 175080 0 0 $X=62680 $Y=174830
X129 36 M4_M3_CDNS_5 $T=62760 191440 0 0 $X=62680 $Y=191190
X130 43 M4_M3_CDNS_5 $T=62760 234970 0 0 $X=62680 $Y=234720
X131 28 M4_M3_CDNS_5 $T=62760 240900 0 0 $X=62680 $Y=240650
X132 7 M4_M3_CDNS_5 $T=62760 242330 0 0 $X=62680 $Y=242080
X133 10 M4_M3_CDNS_5 $T=62760 248290 0 0 $X=62680 $Y=248040
X134 37 M4_M3_CDNS_5 $T=62760 264650 0 0 $X=62680 $Y=264400
X135 23 M4_M3_CDNS_5 $T=62770 81230 0 0 $X=62690 $Y=80980
X136 24 M4_M3_CDNS_5 $T=62770 154450 0 0 $X=62690 $Y=154200
X137 25 M4_M3_CDNS_5 $T=62770 227660 0 0 $X=62690 $Y=227410
X138 41 M4_M3_CDNS_5 $T=63490 16670 0 180 $X=63410 $Y=16420
X139 42 M4_M3_CDNS_5 $T=63490 89890 0 180 $X=63410 $Y=89640
X140 43 M4_M3_CDNS_5 $T=63490 163100 0 180 $X=63410 $Y=162850
X141 38 M4_M3_CDNS_5 $T=63820 12690 0 0 $X=63740 $Y=12440
X142 39 M4_M3_CDNS_5 $T=63820 85910 0 0 $X=63740 $Y=85660
X143 40 M4_M3_CDNS_5 $T=63820 159120 0 0 $X=63740 $Y=158870
X144 11 M4_M3_CDNS_6 $T=11150 139470 0 90 $X=10900 $Y=139390
X145 12 M4_M3_CDNS_6 $T=11150 212690 0 90 $X=10900 $Y=212610
X146 13 M4_M3_CDNS_6 $T=11150 285900 0 90 $X=10900 $Y=285820
X147 14 M4_M3_CDNS_6 $T=16950 140010 0 180 $X=16870 $Y=139760
X148 15 M4_M3_CDNS_6 $T=16950 213230 0 180 $X=16870 $Y=212980
X149 16 M4_M3_CDNS_6 $T=16950 286440 0 180 $X=16870 $Y=286190
X150 20 M4_M3_CDNS_6 $T=31680 139470 0 90 $X=31430 $Y=139390
X151 21 M4_M3_CDNS_6 $T=31680 212690 0 90 $X=31430 $Y=212610
X152 22 M4_M3_CDNS_6 $T=31680 285900 0 90 $X=31430 $Y=285820
X153 17 M4_M3_CDNS_6 $T=41970 139470 0 90 $X=41720 $Y=139390
X154 18 M4_M3_CDNS_6 $T=41970 212690 0 90 $X=41720 $Y=212610
X155 19 M4_M3_CDNS_6 $T=41970 285900 0 90 $X=41720 $Y=285820
X156 29 M4_M3_CDNS_6 $T=51030 71710 0 0 $X=50950 $Y=71460
X157 30 M4_M3_CDNS_6 $T=51030 144930 0 0 $X=50950 $Y=144680
X158 31 M4_M3_CDNS_6 $T=51030 218140 0 0 $X=50950 $Y=217890
X159 35 M4_M3_CDNS_6 $T=51420 72540 0 0 $X=51340 $Y=72290
X160 36 M4_M3_CDNS_6 $T=51420 145760 0 0 $X=51340 $Y=145510
X161 37 M4_M3_CDNS_6 $T=51420 218970 0 0 $X=51340 $Y=218720
X162 32 M4_M3_CDNS_6 $T=54350 80260 0 0 $X=54270 $Y=80010
X163 33 M4_M3_CDNS_6 $T=54350 153480 0 0 $X=54270 $Y=153230
X164 34 M4_M3_CDNS_6 $T=54350 226690 0 0 $X=54270 $Y=226440
X165 26 M4_M3_CDNS_6 $T=63830 19990 0 0 $X=63750 $Y=19740
X166 27 M4_M3_CDNS_6 $T=63830 93210 0 0 $X=63750 $Y=92960
X167 28 M4_M3_CDNS_6 $T=63830 166420 0 0 $X=63750 $Y=166170
X168 2 M5_M4_CDNS_7 $T=49120 82570 0 0 $X=49040 $Y=82320
X169 3 M5_M4_CDNS_7 $T=49120 155790 0 0 $X=49040 $Y=155540
X170 4 M5_M4_CDNS_7 $T=49120 229000 0 0 $X=49040 $Y=228750
X171 23 M5_M4_CDNS_7 $T=53160 72250 0 0 $X=53080 $Y=72000
X172 24 M5_M4_CDNS_7 $T=53160 145470 0 0 $X=53080 $Y=145220
X173 25 M5_M4_CDNS_7 $T=53160 218680 0 0 $X=53080 $Y=218430
X174 23 M5_M4_CDNS_7 $T=55950 72850 0 90 $X=55700 $Y=72770
X175 24 M5_M4_CDNS_7 $T=55950 146070 0 90 $X=55700 $Y=145990
X176 25 M5_M4_CDNS_7 $T=55950 219280 0 90 $X=55700 $Y=219200
X177 2 M5_M4_CDNS_7 $T=62740 103290 0 0 $X=62660 $Y=103040
X178 3 M5_M4_CDNS_7 $T=62740 176510 0 0 $X=62660 $Y=176260
X179 4 M5_M4_CDNS_7 $T=62740 249720 0 0 $X=62660 $Y=249470
X180 38 M5_M4_CDNS_7 $T=62750 87190 0 0 $X=62670 $Y=86940
X181 39 M5_M4_CDNS_7 $T=62750 160410 0 0 $X=62670 $Y=160160
X182 40 M5_M4_CDNS_7 $T=62750 233620 0 0 $X=62670 $Y=233370
X183 41 M5_M4_CDNS_7 $T=62760 88540 0 0 $X=62680 $Y=88290
X184 26 M5_M4_CDNS_7 $T=62760 94470 0 0 $X=62680 $Y=94220
X185 5 M5_M4_CDNS_7 $T=62760 95900 0 0 $X=62680 $Y=95650
X186 8 M5_M4_CDNS_7 $T=62760 101860 0 0 $X=62680 $Y=101610
X187 42 M5_M4_CDNS_7 $T=62760 161760 0 0 $X=62680 $Y=161510
X188 27 M5_M4_CDNS_7 $T=62760 167690 0 0 $X=62680 $Y=167440
X189 6 M5_M4_CDNS_7 $T=62760 169120 0 0 $X=62680 $Y=168870
X190 9 M5_M4_CDNS_7 $T=62760 175080 0 0 $X=62680 $Y=174830
X191 43 M5_M4_CDNS_7 $T=62760 234970 0 0 $X=62680 $Y=234720
X192 28 M5_M4_CDNS_7 $T=62760 240900 0 0 $X=62680 $Y=240650
X193 7 M5_M4_CDNS_7 $T=62760 242330 0 0 $X=62680 $Y=242080
X194 10 M5_M4_CDNS_7 $T=62760 248290 0 0 $X=62680 $Y=248040
X195 23 M5_M4_CDNS_7 $T=62770 81230 0 0 $X=62690 $Y=80980
X196 24 M5_M4_CDNS_7 $T=62770 154450 0 0 $X=62690 $Y=154200
X197 25 M5_M4_CDNS_7 $T=62770 227660 0 0 $X=62690 $Y=227410
X198 41 M5_M4_CDNS_7 $T=63490 16670 0 180 $X=63410 $Y=16420
X199 42 M5_M4_CDNS_7 $T=63490 89890 0 180 $X=63410 $Y=89640
X200 43 M5_M4_CDNS_7 $T=63490 163100 0 180 $X=63410 $Y=162850
X201 38 M5_M4_CDNS_7 $T=63820 12690 0 0 $X=63740 $Y=12440
X202 39 M5_M4_CDNS_7 $T=63820 85910 0 0 $X=63740 $Y=85660
X203 40 M5_M4_CDNS_7 $T=63820 159120 0 0 $X=63740 $Y=158870
X204 8 M4_M3_CDNS_8 $T=50440 71360 0 0 $X=50360 $Y=71230
X205 9 M4_M3_CDNS_8 $T=50440 144580 0 0 $X=50360 $Y=144450
X206 10 M4_M3_CDNS_8 $T=50440 217790 0 0 $X=50360 $Y=217660
X207 5 M4_M3_CDNS_8 $T=50730 70270 0 90 $X=50600 $Y=70190
X208 6 M4_M3_CDNS_8 $T=50730 143490 0 90 $X=50600 $Y=143410
X209 7 M4_M3_CDNS_8 $T=50730 216700 0 90 $X=50600 $Y=216620
X210 2 M4_M3_CDNS_8 $T=57550 91880 0 0 $X=57470 $Y=91750
X211 3 M4_M3_CDNS_8 $T=57550 165100 0 0 $X=57470 $Y=164970
X212 4 M4_M3_CDNS_8 $T=57550 238310 0 0 $X=57470 $Y=238180
X213 23 M4_M3_CDNS_8 $T=63870 9350 0 0 $X=63790 $Y=9220
X214 24 M4_M3_CDNS_8 $T=63870 82570 0 0 $X=63790 $Y=82440
X215 25 M4_M3_CDNS_8 $T=63870 155780 0 0 $X=63790 $Y=155650
X216 4 M3_M2_CDNS_9 $T=62210 216190 0 90 $X=61960 $Y=216110
X217 3 M3_M2_CDNS_9 $T=62240 142980 0 90 $X=61990 $Y=142900
X218 2 M3_M2_CDNS_9 $T=62300 69760 0 90 $X=62050 $Y=69680
X219 32 M3_M2_CDNS_9 $T=62650 125410 0 0 $X=62570 $Y=125160
X220 33 M3_M2_CDNS_9 $T=62650 198630 0 0 $X=62570 $Y=198380
X221 2 M3_M2_CDNS_9 $T=62740 103290 0 0 $X=62660 $Y=103040
X222 3 M3_M2_CDNS_9 $T=62740 176510 0 0 $X=62660 $Y=176260
X223 4 M3_M2_CDNS_9 $T=62740 249720 0 0 $X=62660 $Y=249470
X224 34 M3_M2_CDNS_9 $T=62740 271840 0 0 $X=62660 $Y=271590
X225 38 M3_M2_CDNS_9 $T=62750 87190 0 0 $X=62670 $Y=86940
X226 29 M3_M2_CDNS_9 $T=62750 111060 0 0 $X=62670 $Y=110810
X227 39 M3_M2_CDNS_9 $T=62750 160410 0 0 $X=62670 $Y=160160
X228 30 M3_M2_CDNS_9 $T=62750 184280 0 0 $X=62670 $Y=184030
X229 40 M3_M2_CDNS_9 $T=62750 233620 0 0 $X=62670 $Y=233370
X230 31 M3_M2_CDNS_9 $T=62750 257490 0 0 $X=62670 $Y=257240
X231 41 M3_M2_CDNS_9 $T=62760 88540 0 0 $X=62680 $Y=88290
X232 26 M3_M2_CDNS_9 $T=62760 94470 0 0 $X=62680 $Y=94220
X233 5 M3_M2_CDNS_9 $T=62760 95900 0 0 $X=62680 $Y=95650
X234 8 M3_M2_CDNS_9 $T=62760 101860 0 0 $X=62680 $Y=101610
X235 35 M3_M2_CDNS_9 $T=62760 118220 0 0 $X=62680 $Y=117970
X236 42 M3_M2_CDNS_9 $T=62760 161760 0 0 $X=62680 $Y=161510
X237 27 M3_M2_CDNS_9 $T=62760 167690 0 0 $X=62680 $Y=167440
X238 6 M3_M2_CDNS_9 $T=62760 169120 0 0 $X=62680 $Y=168870
X239 9 M3_M2_CDNS_9 $T=62760 175080 0 0 $X=62680 $Y=174830
X240 36 M3_M2_CDNS_9 $T=62760 191440 0 0 $X=62680 $Y=191190
X241 43 M3_M2_CDNS_9 $T=62760 234970 0 0 $X=62680 $Y=234720
X242 28 M3_M2_CDNS_9 $T=62760 240900 0 0 $X=62680 $Y=240650
X243 7 M3_M2_CDNS_9 $T=62760 242330 0 0 $X=62680 $Y=242080
X244 10 M3_M2_CDNS_9 $T=62760 248290 0 0 $X=62680 $Y=248040
X245 37 M3_M2_CDNS_9 $T=62760 264650 0 0 $X=62680 $Y=264400
X246 23 M3_M2_CDNS_9 $T=62770 81230 0 0 $X=62690 $Y=80980
X247 24 M3_M2_CDNS_9 $T=62770 154450 0 0 $X=62690 $Y=154200
X248 25 M3_M2_CDNS_9 $T=62770 227660 0 0 $X=62690 $Y=227410
X249 41 M3_M2_CDNS_9 $T=63490 16670 0 180 $X=63410 $Y=16420
X250 42 M3_M2_CDNS_9 $T=63490 89890 0 180 $X=63410 $Y=89640
X251 43 M3_M2_CDNS_9 $T=63490 163100 0 180 $X=63410 $Y=162850
X252 38 M3_M2_CDNS_9 $T=63820 12690 0 0 $X=63740 $Y=12440
X253 39 M3_M2_CDNS_9 $T=63820 85910 0 0 $X=63740 $Y=85660
X254 40 M3_M2_CDNS_9 $T=63820 159120 0 0 $X=63740 $Y=158870
X255 26 M3_M2_CDNS_9 $T=63830 19990 0 0 $X=63750 $Y=19740
X256 27 M3_M2_CDNS_9 $T=63830 93210 0 0 $X=63750 $Y=92960
X257 28 M3_M2_CDNS_9 $T=63830 166420 0 0 $X=63750 $Y=166170
X258 23 M3_M2_CDNS_9 $T=63870 9350 0 0 $X=63790 $Y=9100
X259 24 M3_M2_CDNS_9 $T=63870 82570 0 0 $X=63790 $Y=82320
X260 25 M3_M2_CDNS_9 $T=63870 155780 0 0 $X=63790 $Y=155530
X261 4 M2_M1_CDNS_10 $T=62210 216190 0 90 $X=61960 $Y=216110
X262 3 M2_M1_CDNS_10 $T=62240 142980 0 90 $X=61990 $Y=142900
X263 2 M2_M1_CDNS_10 $T=62300 69760 0 90 $X=62050 $Y=69680
X264 32 M2_M1_CDNS_10 $T=62650 125410 0 0 $X=62570 $Y=125160
X265 33 M2_M1_CDNS_10 $T=62650 198630 0 0 $X=62570 $Y=198380
X266 2 M2_M1_CDNS_10 $T=62740 103290 0 0 $X=62660 $Y=103040
X267 3 M2_M1_CDNS_10 $T=62740 176510 0 0 $X=62660 $Y=176260
X268 4 M2_M1_CDNS_10 $T=62740 249720 0 0 $X=62660 $Y=249470
X269 34 M2_M1_CDNS_10 $T=62740 271840 0 0 $X=62660 $Y=271590
X270 38 M2_M1_CDNS_10 $T=62750 87190 0 0 $X=62670 $Y=86940
X271 29 M2_M1_CDNS_10 $T=62750 111060 0 0 $X=62670 $Y=110810
X272 39 M2_M1_CDNS_10 $T=62750 160410 0 0 $X=62670 $Y=160160
X273 30 M2_M1_CDNS_10 $T=62750 184280 0 0 $X=62670 $Y=184030
X274 40 M2_M1_CDNS_10 $T=62750 233620 0 0 $X=62670 $Y=233370
X275 31 M2_M1_CDNS_10 $T=62750 257490 0 0 $X=62670 $Y=257240
X276 41 M2_M1_CDNS_10 $T=62760 88540 0 0 $X=62680 $Y=88290
X277 26 M2_M1_CDNS_10 $T=62760 94470 0 0 $X=62680 $Y=94220
X278 5 M2_M1_CDNS_10 $T=62760 95900 0 0 $X=62680 $Y=95650
X279 8 M2_M1_CDNS_10 $T=62760 101860 0 0 $X=62680 $Y=101610
X280 35 M2_M1_CDNS_10 $T=62760 118220 0 0 $X=62680 $Y=117970
X281 42 M2_M1_CDNS_10 $T=62760 161760 0 0 $X=62680 $Y=161510
X282 27 M2_M1_CDNS_10 $T=62760 167690 0 0 $X=62680 $Y=167440
X283 6 M2_M1_CDNS_10 $T=62760 169120 0 0 $X=62680 $Y=168870
X284 9 M2_M1_CDNS_10 $T=62760 175080 0 0 $X=62680 $Y=174830
X285 36 M2_M1_CDNS_10 $T=62760 191440 0 0 $X=62680 $Y=191190
X286 43 M2_M1_CDNS_10 $T=62760 234970 0 0 $X=62680 $Y=234720
X287 28 M2_M1_CDNS_10 $T=62760 240900 0 0 $X=62680 $Y=240650
X288 7 M2_M1_CDNS_10 $T=62760 242330 0 0 $X=62680 $Y=242080
X289 10 M2_M1_CDNS_10 $T=62760 248290 0 0 $X=62680 $Y=248040
X290 37 M2_M1_CDNS_10 $T=62760 264650 0 0 $X=62680 $Y=264400
X291 23 M2_M1_CDNS_10 $T=62770 81230 0 0 $X=62690 $Y=80980
X292 24 M2_M1_CDNS_10 $T=62770 154450 0 0 $X=62690 $Y=154200
X293 25 M2_M1_CDNS_10 $T=62770 227660 0 0 $X=62690 $Y=227410
X294 41 M2_M1_CDNS_10 $T=63490 16670 0 180 $X=63410 $Y=16420
X295 42 M2_M1_CDNS_10 $T=63490 89890 0 180 $X=63410 $Y=89640
X296 43 M2_M1_CDNS_10 $T=63490 163100 0 180 $X=63410 $Y=162850
X297 38 M2_M1_CDNS_10 $T=63820 12690 0 0 $X=63740 $Y=12440
X298 39 M2_M1_CDNS_10 $T=63820 85910 0 0 $X=63740 $Y=85660
X299 40 M2_M1_CDNS_10 $T=63820 159120 0 0 $X=63740 $Y=158870
X300 26 M2_M1_CDNS_10 $T=63830 19990 0 0 $X=63750 $Y=19740
X301 27 M2_M1_CDNS_10 $T=63830 93210 0 0 $X=63750 $Y=92960
X302 28 M2_M1_CDNS_10 $T=63830 166420 0 0 $X=63750 $Y=166170
X303 23 M2_M1_CDNS_10 $T=63870 9350 0 0 $X=63790 $Y=9100
X304 24 M2_M1_CDNS_10 $T=63870 82570 0 0 $X=63790 $Y=82320
X305 25 M2_M1_CDNS_10 $T=63870 155780 0 0 $X=63790 $Y=155530
X306 32 M2_M1_CDNS_11 $T=63810 53250 0 0 $X=63730 $Y=53120
X307 33 M2_M1_CDNS_11 $T=63810 126470 0 0 $X=63730 $Y=126340
X308 34 M2_M1_CDNS_11 $T=63810 199680 0 0 $X=63730 $Y=199550
X309 35 M2_M1_CDNS_11 $T=63830 45950 0 0 $X=63750 $Y=45820
X310 36 M2_M1_CDNS_11 $T=63830 119170 0 0 $X=63750 $Y=119040
X311 37 M2_M1_CDNS_11 $T=63830 192380 0 0 $X=63750 $Y=192250
X312 29 M2_M1_CDNS_11 $T=63860 38630 0 0 $X=63780 $Y=38500
X313 30 M2_M1_CDNS_11 $T=63860 111850 0 0 $X=63780 $Y=111720
X314 31 M2_M1_CDNS_11 $T=63860 185060 0 0 $X=63780 $Y=184930
X315 2 M4_M3_CDNS_12 $T=49120 82570 0 0 $X=49040 $Y=82320
X316 3 M4_M3_CDNS_12 $T=49120 155790 0 0 $X=49040 $Y=155540
X317 4 M4_M3_CDNS_12 $T=49120 229000 0 0 $X=49040 $Y=228750
X318 23 M4_M3_CDNS_12 $T=53160 72250 0 0 $X=53080 $Y=72000
X319 24 M4_M3_CDNS_12 $T=53160 145470 0 0 $X=53080 $Y=145220
X320 25 M4_M3_CDNS_12 $T=53160 218680 0 0 $X=53080 $Y=218430
X321 23 M4_M3_CDNS_12 $T=55950 72850 0 90 $X=55700 $Y=72770
X322 24 M4_M3_CDNS_12 $T=55950 146070 0 90 $X=55700 $Y=145990
X323 25 M4_M3_CDNS_12 $T=55950 219280 0 90 $X=55700 $Y=219200
X324 44 11 20 17 45 1 46 47 48 14
+ 49 50 51 52 53 54 55 56 57 58
+ 59 60 61 62 63 41 32 2 38 35
+ 26 5 29 23 8 64 65 66 67 68
+ 69 70 71 72 73 221 1391 1412 162 220
+ 217 167 356 163 161 135 166 242 1340 1393
+ 1395 218 216 164 1394 1423 1390 219 192 1392
+ 165 1455 1396 1450 2167 2103 2104 2105 2106 2170
+ 144 153 178 186 187 193 223 224 257 259
+ 271 273 276 299 314 315 2172 2107 2108 2109
+ 2110 2174 2175 2111 2112 2113 2114 2178 2180 2115
+ 2116 2117 2118 2182 2169 2173 2177 2181 2168 2171
+ 2176 2179 ph2p2_processing_element $T=370 -60 0 0 $X=260 $Y=-60
X325 74 12 21 18 45 1 46 75 48 15
+ 76 11 77 78 79 14 80 81 82 20
+ 83 84 17 85 86 42 33 3 39 36
+ 27 6 30 24 9 23 38 41 26 5
+ 8 2 29 35 32 513 1593 1614 454 512
+ 509 459 648 455 453 427 458 534 1542 1595
+ 1597 510 508 456 1596 1625 1592 511 484 1594
+ 457 1657 1598 1652 2183 2119 2120 2121 2122 2186
+ 436 445 470 478 479 485 515 516 549 551
+ 563 565 568 591 606 607 2188 2123 2124 2125
+ 2126 2190 2191 2127 2128 2129 2130 2194 2196 2131
+ 2132 2133 2134 2198 2185 2189 2193 2197 2184 2187
+ 2192 2195 ph2p2_processing_element $T=370 73140 0 0 $X=260 $Y=73140
X326 87 13 22 19 45 1 46 88 48 16
+ 89 12 90 91 92 15 93 94 95 21
+ 96 97 18 98 99 43 34 4 40 37
+ 28 7 31 25 10 24 39 42 27 6
+ 9 3 30 36 33 805 1795 1816 746 804
+ 801 751 940 747 745 719 750 826 1744 1797
+ 1799 802 800 748 1798 1827 1794 803 776 1796
+ 749 1859 1800 1854 2199 2135 2136 2137 2138 2202
+ 728 737 762 770 771 777 807 808 841 843
+ 855 857 860 883 898 899 2204 2139 2140 2141
+ 2142 2206 2207 2143 2144 2145 2146 2210 2212 2147
+ 2148 2149 2150 2214 2201 2205 2209 2213 2200 2203
+ 2208 2211 ph2p2_processing_element $T=370 146340 0 0 $X=260 $Y=146340
X327 100 101 102 103 45 1 46 104 48 105
+ 106 13 107 108 109 16 110 111 112 22
+ 113 114 19 115 116 117 118 119 120 121
+ 122 123 124 125 126 25 40 43 28 7
+ 10 4 31 37 34 1097 1997 2018 1038 1096
+ 1093 1043 1232 1039 1037 1011 1042 1118 1946 1999
+ 2001 1094 1092 1040 2000 2029 1996 1095 1068 1998
+ 1041 2061 2002 2056 2215 2151 2152 2153 2154 2218
+ 1020 1029 1054 1062 1063 1069 1099 1100 1133 1135
+ 1147 1149 1152 1175 1190 1191 2220 2155 2156 2157
+ 2158 2222 2223 2159 2160 2161 2162 2226 2228 2163
+ 2164 2165 2166 2230 2217 2221 2225 2229 2216 2219
+ 2224 2227 ph2p2_processing_element $T=370 219540 0 0 $X=260 $Y=219540
M0 2106 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=72010 $dt=1
M1 2122 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=145210 $dt=1
M2 2138 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=218410 $dt=1
M3 2154 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=2290 $Y=291610 $dt=1
M4 153 135 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.8911 scb=0.00996238 scc=0.000256798 $X=2380 $Y=920 $dt=1
M5 445 427 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=74120 $dt=1
M6 737 719 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=147320 $dt=1
M7 1029 1011 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=220520 $dt=1
M8 2167 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=72040 $dt=1
M9 2183 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=145240 $dt=1
M10 2199 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=218440 $dt=1
M11 2215 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=3620 $Y=291640 $dt=1
M12 2168 135 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=3710 $Y=680 $dt=1
M13 2184 427 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=73880 $dt=1
M14 2200 719 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=147080 $dt=1
M15 2216 1011 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=220280 $dt=1
M16 178 144 2168 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=4680 $Y=620 $dt=1
M17 470 436 2184 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=73820 $dt=1
M18 762 728 2200 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=147020 $dt=1
M19 1054 1020 2216 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=220220 $dt=1
M20 2103 46 11 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=72040 $dt=1
M21 2119 46 12 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=145240 $dt=1
M22 2135 46 13 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=218440 $dt=1
M23 2151 46 101 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=4800 $Y=291640 $dt=1
M24 178 153 2168 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=5640 $Y=620 $dt=1
M25 470 445 2184 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=73820 $dt=1
M26 762 737 2200 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=147020 $dt=1
M27 1054 1029 2216 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=220220 $dt=1
M28 2105 2103 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=71950 $dt=1
M29 2121 2119 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=145150 $dt=1
M30 2137 2135 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=218350 $dt=1
M31 2153 2151 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=6000 $Y=291550 $dt=1
M32 2168 47 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=6600 $Y=620 $dt=1
M33 2184 75 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=73820 $dt=1
M34 2200 88 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=147020 $dt=1
M35 2216 104 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=220220 $dt=1
M36 2105 2104 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=71960 $dt=1
M37 2121 2120 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=145160 $dt=1
M38 2137 2136 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=218360 $dt=1
M39 2153 2152 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=7240 $Y=291560 $dt=1
M40 186 193 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=8260 $Y=920 $dt=1
M41 478 485 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=74120 $dt=1
M42 770 777 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=147320 $dt=1
M43 1062 1069 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=220520 $dt=1
M44 2169 2105 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=72010 $dt=1
M45 2185 2121 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=145210 $dt=1
M46 2201 2137 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=218410 $dt=1
M47 2217 2153 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=8490 $Y=291610 $dt=1
M48 187 178 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=9220 $Y=920 $dt=1
M49 479 470 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=74120 $dt=1
M50 771 762 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=147320 $dt=1
M51 1063 1054 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=220520 $dt=1
M52 2170 2106 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=72040 $dt=1
M53 2186 2122 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=145240 $dt=1
M54 2202 2138 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=218440 $dt=1
M55 2218 2154 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=9820 $Y=291640 $dt=1
M56 2171 178 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=10550 $Y=680 $dt=1
M57 2187 470 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=73880 $dt=1
M58 2203 762 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=147080 $dt=1
M59 2219 1054 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=220280 $dt=1
M60 2103 2106 2169 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=72040 $dt=1
M61 2119 2122 2185 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=145240 $dt=1
M62 2135 2138 2201 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=218440 $dt=1
M63 2151 2154 2217 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=11000 $Y=291640 $dt=1
M64 1340 186 2171 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=11520 $Y=620 $dt=1
M65 1542 478 2187 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=73820 $dt=1
M66 1744 770 2203 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=147020 $dt=1
M67 1946 1062 2219 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=220220 $dt=1
M68 1340 187 2171 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=12480 $Y=620 $dt=1
M69 1542 479 2187 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=73820 $dt=1
M70 1744 771 2203 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=147020 $dt=1
M71 1946 1063 2219 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=220220 $dt=1
M72 2110 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=72010 $dt=1
M73 2126 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=145210 $dt=1
M74 2142 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=218410 $dt=1
M75 2158 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=12530 $Y=291610 $dt=1
M76 2171 193 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=13440 $Y=620 $dt=1
M77 2187 485 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=73820 $dt=1
M78 2203 777 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=147020 $dt=1
M79 2219 1069 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=220220 $dt=1
M80 2172 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=72040 $dt=1
M81 2188 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=145240 $dt=1
M82 2204 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=218440 $dt=1
M83 2220 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=13860 $Y=291640 $dt=1
M84 2107 46 14 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=72040 $dt=1
M85 2123 46 15 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=145240 $dt=1
M86 2139 46 16 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=218440 $dt=1
M87 2155 46 105 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=15040 $Y=291640 $dt=1
M88 223 193 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=15510 $Y=650 $dt=1
M89 515 485 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=73850 $dt=1
M90 807 777 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=147050 $dt=1
M91 1099 1069 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=220250 $dt=1
M92 48 178 223 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=15920 $Y=650 $dt=1
M93 48 470 515 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=73850 $dt=1
M94 48 762 807 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=147050 $dt=1
M95 48 1054 1099 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=220250 $dt=1
M96 2109 2107 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=71950 $dt=1
M97 2125 2123 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=145150 $dt=1
M98 2141 2139 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=218350 $dt=1
M99 2157 2155 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=16240 $Y=291550 $dt=1
M100 2109 2108 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=71960 $dt=1
M101 2125 2124 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=145160 $dt=1
M102 2141 2140 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=218360 $dt=1
M103 2157 2156 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=17480 $Y=291560 $dt=1
M104 224 47 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=18490 $Y=910 $dt=1
M105 516 75 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=74110 $dt=1
M106 808 88 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=147310 $dt=1
M107 1100 104 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=220510 $dt=1
M108 2173 2109 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=72010 $dt=1
M109 2189 2125 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=145210 $dt=1
M110 2205 2141 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=218410 $dt=1
M111 2221 2157 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=18730 $Y=291610 $dt=1
M112 48 135 224 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=18900 $Y=910 $dt=1
M113 48 427 516 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=74110 $dt=1
M114 48 719 808 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=147310 $dt=1
M115 48 1011 1100 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=220510 $dt=1
M116 2174 2110 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=72040 $dt=1
M117 2190 2126 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=145240 $dt=1
M118 2206 2142 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=218440 $dt=1
M119 2222 2158 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=20060 $Y=291640 $dt=1
M120 2107 2110 2173 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=72040 $dt=1
M121 2123 2126 2189 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=145240 $dt=1
M122 2139 2142 2205 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=218440 $dt=1
M123 2155 2158 2221 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=21240 $Y=291640 $dt=1
M124 299 223 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=21330 $Y=910 $dt=1
M125 591 515 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=74110 $dt=1
M126 883 807 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=147310 $dt=1
M127 1175 1099 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=220510 $dt=1
M128 48 224 299 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=21740 $Y=910 $dt=1
M129 48 516 591 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=74110 $dt=1
M130 48 808 883 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=147310 $dt=1
M131 48 1100 1175 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=220510 $dt=1
M132 2114 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=72010 $dt=1
M133 2130 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=145210 $dt=1
M134 2146 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=218410 $dt=1
M135 2162 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=22770 $Y=291610 $dt=1
M136 257 56 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=23380 $Y=920 $dt=1
M137 549 81 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=74120 $dt=1
M138 841 94 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=147320 $dt=1
M139 1133 111 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=220520 $dt=1
M140 2175 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=72040 $dt=1
M141 2191 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=145240 $dt=1
M142 2207 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=218440 $dt=1
M143 2223 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=24100 $Y=291640 $dt=1
M144 259 242 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=24340 $Y=920 $dt=1
M145 551 534 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=74120 $dt=1
M146 843 826 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=147320 $dt=1
M147 1135 1118 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=220520 $dt=1
M148 2111 46 20 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=72040 $dt=1
M149 2127 46 21 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=145240 $dt=1
M150 2143 46 22 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=218440 $dt=1
M151 2159 46 102 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=25280 $Y=291640 $dt=1
M152 2176 242 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=25670 $Y=680 $dt=1
M153 2192 534 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=73880 $dt=1
M154 2208 826 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=147080 $dt=1
M155 2224 1118 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=220280 $dt=1
M156 2113 2111 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=71950 $dt=1
M157 2129 2127 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=145150 $dt=1
M158 2145 2143 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=218350 $dt=1
M159 2161 2159 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=26480 $Y=291550 $dt=1
M160 271 257 2176 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=26640 $Y=620 $dt=1
M161 563 549 2192 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=73820 $dt=1
M162 855 841 2208 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=147020 $dt=1
M163 1147 1133 2224 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=220220 $dt=1
M164 271 259 2176 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=27600 $Y=620 $dt=1
M165 563 551 2192 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=73820 $dt=1
M166 855 843 2208 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=147020 $dt=1
M167 1147 1135 2224 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=220220 $dt=1
M168 2113 2112 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=71960 $dt=1
M169 2129 2128 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=145160 $dt=1
M170 2145 2144 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=218360 $dt=1
M171 2161 2160 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=27720 $Y=291560 $dt=1
M172 2176 56 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=28560 $Y=620 $dt=1
M173 2192 81 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=73820 $dt=1
M174 2208 94 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=147020 $dt=1
M175 2224 111 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=220220 $dt=1
M176 2177 2113 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=72010 $dt=1
M177 2193 2129 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=145210 $dt=1
M178 2209 2145 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=218410 $dt=1
M179 2225 2161 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=28970 $Y=291610 $dt=1
M180 273 299 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=30220 $Y=920 $dt=1
M181 565 591 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=74120 $dt=1
M182 857 883 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=147320 $dt=1
M183 1149 1175 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=220520 $dt=1
M184 2178 2114 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=72040 $dt=1
M185 2194 2130 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=145240 $dt=1
M186 2210 2146 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=218440 $dt=1
M187 2226 2162 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=30300 $Y=291640 $dt=1
M188 276 271 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=31180 $Y=920 $dt=1
M189 568 563 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=74120 $dt=1
M190 860 855 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=147320 $dt=1
M191 1152 1147 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=220520 $dt=1
M192 2111 2114 2177 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=72040 $dt=1
M193 2127 2130 2193 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=145240 $dt=1
M194 2143 2146 2209 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=218440 $dt=1
M195 2159 2162 2225 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=31480 $Y=291640 $dt=1
M196 2179 271 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=32510 $Y=680 $dt=1
M197 2195 563 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=73880 $dt=1
M198 2211 855 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=147080 $dt=1
M199 2227 1147 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=220280 $dt=1
M200 2118 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=72010 $dt=1
M201 2134 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=145210 $dt=1
M202 2150 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=218410 $dt=1
M203 2166 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=33010 $Y=291610 $dt=1
M204 1423 273 2179 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=33480 $Y=620 $dt=1
M205 1625 565 2195 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=73820 $dt=1
M206 1827 857 2211 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=147020 $dt=1
M207 2029 1149 2227 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=220220 $dt=1
M208 2180 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=72040 $dt=1
M209 2196 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=145240 $dt=1
M210 2212 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=218440 $dt=1
M211 2228 46 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=34340 $Y=291640 $dt=1
M212 1423 276 2179 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=34440 $Y=620 $dt=1
M213 1625 568 2195 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=73820 $dt=1
M214 1827 860 2211 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=147020 $dt=1
M215 2029 1152 2227 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=220220 $dt=1
M216 2179 299 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=35400 $Y=620 $dt=1
M217 2195 591 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=73820 $dt=1
M218 2211 883 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=147020 $dt=1
M219 2227 1175 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=220220 $dt=1
M220 2115 46 17 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=72040 $dt=1
M221 2131 46 18 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=145240 $dt=1
M222 2147 46 19 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=218440 $dt=1
M223 2163 46 103 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=35520 $Y=291640 $dt=1
M224 2117 2115 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=71950 $dt=1
M225 2133 2131 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=145150 $dt=1
M226 2149 2147 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=218350 $dt=1
M227 2165 2163 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=36720 $Y=291550 $dt=1
M228 314 299 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=37470 $Y=650 $dt=1
M229 606 591 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=73850 $dt=1
M230 898 883 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=147050 $dt=1
M231 1190 1175 48 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=220250 $dt=1
M232 48 271 314 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=37880 $Y=650 $dt=1
M233 48 563 606 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=73850 $dt=1
M234 48 855 898 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=147050 $dt=1
M235 48 1147 1190 48 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=220250 $dt=1
M236 2117 2116 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=71960 $dt=1
M237 2133 2132 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=145160 $dt=1
M238 2149 2148 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=218360 $dt=1
M239 2165 2164 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=37960 $Y=291560 $dt=1
M240 2181 2117 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=72010 $dt=1
M241 2197 2133 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=145210 $dt=1
M242 2213 2149 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=218410 $dt=1
M243 2229 2165 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=39210 $Y=291610 $dt=1
M244 315 56 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=40450 $Y=910 $dt=1
M245 607 81 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=74110 $dt=1
M246 899 94 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=147310 $dt=1
M247 1191 111 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=220510 $dt=1
M248 2182 2118 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=72040 $dt=1
M249 2198 2134 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=145240 $dt=1
M250 2214 2150 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=218440 $dt=1
M251 2230 2166 48 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=40540 $Y=291640 $dt=1
M252 48 242 315 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=40860 $Y=910 $dt=1
M253 48 534 607 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=74110 $dt=1
M254 48 826 899 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=147310 $dt=1
M255 48 1118 1191 48 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=220510 $dt=1
M256 2115 2118 2181 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=72040 $dt=1
M257 2131 2134 2197 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=145240 $dt=1
M258 2147 2150 2213 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=218440 $dt=1
M259 2163 2166 2229 48 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=41720 $Y=291640 $dt=1
.ends ph2p3_Matrix_vector_Multiplication
