* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 1_bit_Full_Adder_ver2                        *
* Netlisted  : Wed Oct 16 07:19:28 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_9                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_9 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_10                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_10 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR2_1X                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR2_1X 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=10
X0 6 M2_M1_CDNS_6 $T=1040 1920 0 90 $X=910 $Y=1840
X1 7 M2_M1_CDNS_6 $T=1960 1580 0 90 $X=1830 $Y=1500
X2 8 M2_M1_CDNS_6 $T=3270 3070 0 0 $X=3190 $Y=2940
X3 9 M2_M1_CDNS_6 $T=3360 690 0 90 $X=3230 $Y=610
X4 6 M2_M1_CDNS_6 $T=3460 1920 0 90 $X=3330 $Y=1840
X5 8 M2_M1_CDNS_6 $T=3790 3050 0 0 $X=3710 $Y=2920
X6 7 M2_M1_CDNS_6 $T=4520 1580 0 90 $X=4390 $Y=1500
X7 8 M2_M1_CDNS_6 $T=4720 3050 0 0 $X=4640 $Y=2920
X8 9 M2_M1_CDNS_6 $T=5550 690 0 90 $X=5420 $Y=610
X9 8 M2_M1_CDNS_6 $T=5650 3050 0 0 $X=5570 $Y=2920
X10 1 M1_PO_CDNS_7 $T=580 2010 0 90 $X=460 $Y=1910
X11 2 M1_PO_CDNS_7 $T=1490 1580 0 90 $X=1370 $Y=1480
X12 6 M1_PO_CDNS_7 $T=3880 1920 0 90 $X=3760 $Y=1820
X13 7 M1_PO_CDNS_7 $T=4800 1580 0 90 $X=4680 $Y=1480
X14 4 1 6 4 nmos1v_CDNS_9 $T=650 860 0 0 $X=230 $Y=660
X15 4 2 7 4 nmos1v_CDNS_9 $T=1580 860 0 0 $X=1160 $Y=660
X16 4 2 9 4 nmos1v_CDNS_9 $T=3020 860 0 0 $X=2600 $Y=660
X17 10 6 5 4 nmos1v_CDNS_9 $T=3950 860 0 0 $X=3530 $Y=660
X18 10 7 4 4 nmos1v_CDNS_9 $T=4880 860 0 0 $X=4460 $Y=660
X19 9 1 5 4 nmos1v_CDNS_9 $T=5810 860 0 0 $X=5390 $Y=660
X20 3 6 1 4 3 pmos1v_CDNS_10 $T=650 2490 0 0 $X=230 $Y=2290
X21 3 7 2 4 3 pmos1v_CDNS_10 $T=1580 2490 0 0 $X=1160 $Y=2290
X22 3 8 2 4 3 pmos1v_CDNS_10 $T=3020 2500 0 0 $X=2600 $Y=2300
X23 8 5 6 4 3 pmos1v_CDNS_10 $T=3950 2500 0 0 $X=3530 $Y=2300
X24 8 5 7 4 3 pmos1v_CDNS_10 $T=4880 2500 0 0 $X=4460 $Y=2300
X25 8 3 1 4 3 pmos1v_CDNS_10 $T=5810 2500 0 0 $X=5390 $Y=2300
M0 8 2 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3020 $Y=2500 $dt=1
M1 5 6 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3950 $Y=2500 $dt=1
M2 5 7 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=4880 $Y=2500 $dt=1
M3 3 1 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=5810 $Y=2500 $dt=1
.ends XOR2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_13                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_13 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_7 $T=520 1770 0 90 $X=400 $Y=1670
X1 4 M1_PO_CDNS_7 $T=1200 1830 0 90 $X=1080 $Y=1730
X2 2 3 cellTmpl_CDNS_13 $T=120 150 0 0 $X=0 $Y=10
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=620 $Y=720 $dt=0
M1 5 4 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=830 $Y=720 $dt=0
.ends NAND2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X 1 2 3 4
** N=4 EP=4 FDC=2
X0 3 M1_PO_CDNS_7 $T=970 1740 0 90 $X=850 $Y=1640
X1 1 2 cellTmpl_CDNS_13 $T=130 140 0 0 $X=10 $Y=0
M0 4 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6908 scb=0.0179614 scc=0.00130074 $X=1090 $Y=1110 $dt=0
M1 4 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=18.2452 scb=0.0177397 scc=0.00150411 $X=1090 $Y=2120 $dt=1
.ends INV_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 1_bit_Full_Adder_ver2                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 1_bit_Full_Adder_ver2 4 1 2 13 9 7 6
** N=28 EP=7 FDC=46
X0 1 M3_M2_CDNS_1 $T=1190 1430 0 0 $X=1110 $Y=1180
X1 2 M3_M2_CDNS_1 $T=7590 1430 0 0 $X=7510 $Y=1180
X2 1 M3_M2_CDNS_1 $T=14680 1820 0 90 $X=14430 $Y=1740
X3 3 M3_M2_CDNS_1 $T=14880 1070 0 90 $X=14630 $Y=990
X4 2 M3_M2_CDNS_1 $T=16700 1810 0 90 $X=16450 $Y=1730
X5 3 M3_M2_CDNS_1 $T=18700 1820 0 90 $X=18450 $Y=1740
X6 1 M3_M2_CDNS_1 $T=21290 1610 0 180 $X=21210 $Y=1360
X7 2 M3_M2_CDNS_1 $T=22680 1820 0 90 $X=22430 $Y=1740
X8 1 M2_M1_CDNS_2 $T=1190 1430 0 0 $X=1110 $Y=1180
X9 2 M2_M1_CDNS_2 $T=7590 1430 0 0 $X=7510 $Y=1180
X10 1 M2_M1_CDNS_2 $T=14680 1820 0 90 $X=14430 $Y=1740
X11 3 M2_M1_CDNS_2 $T=14880 1070 0 90 $X=14630 $Y=990
X12 2 M2_M1_CDNS_2 $T=16700 1810 0 90 $X=16450 $Y=1730
X13 3 M2_M1_CDNS_2 $T=18700 1820 0 90 $X=18450 $Y=1740
X14 1 M2_M1_CDNS_2 $T=21290 1610 0 180 $X=21210 $Y=1360
X15 2 M2_M1_CDNS_2 $T=22680 1820 0 90 $X=22430 $Y=1740
X16 4 M4_M3_CDNS_3 $T=270 1860 0 0 $X=190 $Y=1610
X17 4 M4_M3_CDNS_3 $T=13290 1610 0 0 $X=13210 $Y=1360
X18 4 M4_M3_CDNS_3 $T=15290 1610 0 0 $X=15210 $Y=1360
X19 5 M4_M3_CDNS_3 $T=20710 2200 0 0 $X=20630 $Y=1950
X20 5 M4_M3_CDNS_3 $T=24700 1820 0 90 $X=24450 $Y=1740
X21 4 M3_M2_CDNS_4 $T=270 1860 0 0 $X=190 $Y=1610
X22 4 M3_M2_CDNS_4 $T=13290 1610 0 0 $X=13210 $Y=1360
X23 4 M3_M2_CDNS_4 $T=15290 1610 0 0 $X=15210 $Y=1360
X24 5 M3_M2_CDNS_4 $T=20710 2200 0 0 $X=20630 $Y=1950
X25 5 M3_M2_CDNS_4 $T=24700 1820 0 90 $X=24450 $Y=1740
X26 4 M2_M1_CDNS_5 $T=270 1860 0 0 $X=190 $Y=1610
X27 4 M2_M1_CDNS_5 $T=13290 1610 0 0 $X=13210 $Y=1360
X28 4 M2_M1_CDNS_5 $T=15290 1610 0 0 $X=15210 $Y=1360
X29 5 M2_M1_CDNS_5 $T=20710 2200 0 0 $X=20630 $Y=1950
X30 5 M2_M1_CDNS_5 $T=24700 1820 0 90 $X=24450 $Y=1740
X31 4 1 6 7 8 14 15 27 18 19 XOR2_1X $T=0 0 0 0 $X=0 $Y=0
X32 8 2 6 7 9 16 17 28 20 21 XOR2_1X $T=6400 0 0 0 $X=6400 $Y=0
X33 4 6 7 1 3 22 NAND2_1X $T=13040 -10 0 0 $X=13040 $Y=0
X34 4 6 7 2 10 23 NAND2_1X $T=15040 -10 0 0 $X=15040 $Y=0
X35 10 6 7 3 11 24 NAND2_1X $T=17040 -10 0 0 $X=17040 $Y=0
X36 1 6 7 2 12 25 NAND2_1X $T=21040 -10 0 0 $X=21040 $Y=0
X37 12 6 7 5 13 26 NAND2_1X $T=23040 -10 0 0 $X=23040 $Y=0
X38 6 7 11 5 INV_1X $T=19030 0 0 0 $X=19040 $Y=0
M0 14 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=17.6861 scb=0.0184591 scc=0.000433664 $X=650 $Y=2490 $dt=1
M1 15 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.886 scb=0.00790338 scc=9.25552e-05 $X=1580 $Y=2490 $dt=1
M2 16 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=7050 $Y=2490 $dt=1
M3 17 2 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=7980 $Y=2490 $dt=1
M4 3 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=13660 $Y=2070 $dt=1
M5 6 1 3 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=14070 $Y=2070 $dt=1
M6 10 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=15660 $Y=2070 $dt=1
M7 6 2 10 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=16070 $Y=2070 $dt=1
M8 11 10 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=17660 $Y=2070 $dt=1
M9 6 3 11 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=18070 $Y=2070 $dt=1
M10 12 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=21660 $Y=2070 $dt=1
M11 6 2 12 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=22070 $Y=2070 $dt=1
M12 13 12 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=22.3336 scb=0.0204967 scc=0.00219492 $X=23660 $Y=2070 $dt=1
M13 6 5 13 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=23.6714 scb=0.021925 scc=0.00220002 $X=24070 $Y=2070 $dt=1
.ends 1_bit_Full_Adder_ver2
