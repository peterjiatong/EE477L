* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : NOR2_1X                                      *
* Netlisted  : Mon Sep 30 18:08:53 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_3 D_drain_1 2 3
** N=3 EP=3 FDC=1
M0 D_drain_1 2 3 D_drain_1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.92e-14 PD=5.2e-07 PS=5.6e-07 fw=1.2e-07 sa=3.45e-07 sb=1.4e-07 sca=7.03506 scb=0.00388147 scc=3.26493e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_4 D_drain_1 2 3 B
** N=5 EP=4 FDC=1
M0 D_drain_1 2 3 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=14.9854 scb=0.0121279 scc=0.000129795 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_5                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_5 S_source_0 2 3 B
** N=5 EP=4 FDC=1
M0 3 2 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=15.74 scb=0.0137362 scc=0.000169656 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_6                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_6 D_drain_1 S_source_0 3
** N=3 EP=3 FDC=1
M0 D_drain_1 3 S_source_0 S_source_0 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.92e-14 AS=1.68e-14 PD=5.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=3.45e-07 sca=7.03506 scb=0.00388147 scc=3.26493e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NOR2_1X                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NOR2_1X gnd! in_a in_b out vdd!
** N=6 EP=5 FDC=4
X2 gnd! in_a out nmos1v_CDNS_3 $T=1280 680 0 0 $X=1040 $Y=480
X3 vdd! in_a 6 vdd! pmos1v_CDNS_4 $T=1080 2450 0 0 $X=880 $Y=2250
X4 out in_b 6 vdd! pmos1v_CDNS_5 $T=870 2450 0 0 $X=450 $Y=2250
X5 out gnd! in_b nmos1v_CDNS_6 $T=870 680 0 0 $X=450 $Y=480
.ends NOR2_1X
