* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 1_bit_Full_Adder_ver1                        *
* Netlisted  : Wed Oct 16 05:23:11 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_9                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_9 1 2 3 4 5 6
*.DEVICECLIMB
** N=14 EP=6 FDC=2
M0 4 6 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=500 $Y=570 $dt=0
M1 5 3 4 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=710 $Y=570 $dt=0
.ends cellTmpl_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X 1 2 3 4 5 6
** N=6 EP=6 FDC=4
X0 3 M1_PO_CDNS_6 $T=520 1770 0 90 $X=400 $Y=1670
X1 4 M1_PO_CDNS_6 $T=1200 1830 0 90 $X=1080 $Y=1730
X2 1 2 4 6 5 3 cellTmpl_CDNS_9 $T=120 150 0 0 $X=0 $Y=10
M0 5 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=620 $Y=2080 $dt=1
M1 1 4 5 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=1030 $Y=2080 $dt=1
.ends NAND2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_2X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_2X 1 2 3 4 5 6
** N=6 EP=6 FDC=4
X0 3 M1_PO_CDNS_6 $T=520 1760 0 90 $X=400 $Y=1660
X1 4 M1_PO_CDNS_6 $T=1200 1820 0 90 $X=1080 $Y=1720
X2 1 2 4 6 5 3 cellTmpl_CDNS_9 $T=120 140 0 0 $X=0 $Y=0
M0 5 3 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=15.9511 scb=0.0138709 scc=0.00113792 $X=620 $Y=2070 $dt=1
M1 1 4 5 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=15.9511 scb=0.0138709 scc=0.00113792 $X=1030 $Y=2070 $dt=1
.ends NAND2_2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_14                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_14 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_16                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_16 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_17                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_17 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR2_1X                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR2_1X 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=8
X0 1 M1_PO_CDNS_6 $T=580 2010 0 90 $X=460 $Y=1910
X1 2 M1_PO_CDNS_6 $T=1490 1580 0 90 $X=1370 $Y=1480
X2 6 M1_PO_CDNS_6 $T=3880 1920 0 90 $X=3760 $Y=1820
X3 7 M1_PO_CDNS_6 $T=4800 1580 0 90 $X=4680 $Y=1480
X4 6 M2_M1_CDNS_14 $T=1040 1920 0 90 $X=910 $Y=1840
X5 7 M2_M1_CDNS_14 $T=1960 1580 0 90 $X=1830 $Y=1500
X6 8 M2_M1_CDNS_14 $T=3270 3070 0 0 $X=3190 $Y=2940
X7 9 M2_M1_CDNS_14 $T=3360 690 0 90 $X=3230 $Y=610
X8 6 M2_M1_CDNS_14 $T=3460 1920 0 90 $X=3330 $Y=1840
X9 8 M2_M1_CDNS_14 $T=3790 3050 0 0 $X=3710 $Y=2920
X10 7 M2_M1_CDNS_14 $T=4520 1580 0 90 $X=4390 $Y=1500
X11 8 M2_M1_CDNS_14 $T=4720 3050 0 0 $X=4640 $Y=2920
X12 9 M2_M1_CDNS_14 $T=5550 690 0 90 $X=5420 $Y=610
X13 8 M2_M1_CDNS_14 $T=5650 3050 0 0 $X=5570 $Y=2920
X14 4 1 6 4 nmos1v_CDNS_16 $T=650 860 0 0 $X=230 $Y=660
X15 4 2 7 4 nmos1v_CDNS_16 $T=1580 860 0 0 $X=1160 $Y=660
X16 4 2 9 4 nmos1v_CDNS_16 $T=3020 860 0 0 $X=2600 $Y=660
X17 10 6 5 4 nmos1v_CDNS_16 $T=3950 860 0 0 $X=3530 $Y=660
X18 10 7 4 4 nmos1v_CDNS_16 $T=4880 860 0 0 $X=4460 $Y=660
X19 9 1 5 4 nmos1v_CDNS_16 $T=5810 860 0 0 $X=5390 $Y=660
X20 3 1 6 4 3 pmos1v_CDNS_17 $T=650 2490 0 0 $X=230 $Y=2290
X21 3 2 7 4 3 pmos1v_CDNS_17 $T=1580 2490 0 0 $X=1160 $Y=2290
X22 3 2 8 4 3 pmos1v_CDNS_17 $T=3020 2500 0 0 $X=2600 $Y=2300
X23 8 6 5 4 3 pmos1v_CDNS_17 $T=3950 2500 0 0 $X=3530 $Y=2300
X24 8 7 5 4 3 pmos1v_CDNS_17 $T=4880 2500 0 0 $X=4460 $Y=2300
X25 8 1 3 4 3 pmos1v_CDNS_17 $T=5810 2500 0 0 $X=5390 $Y=2300
M0 8 2 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3020 $Y=2500 $dt=1
M1 5 6 8 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3950 $Y=2500 $dt=1
.ends XOR2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 1_bit_Full_Adder_ver1                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 1_bit_Full_Adder_ver1 4 1 2 3 10 8 7
** N=23 EP=7 FDC=36
X0 1 M3_M2_CDNS_1 $T=1170 1430 0 0 $X=1090 $Y=1180
X1 2 M3_M2_CDNS_1 $T=8020 1830 0 90 $X=7770 $Y=1750
X2 1 M3_M2_CDNS_1 $T=8650 1560 0 0 $X=8570 $Y=1310
X3 3 M3_M2_CDNS_1 $T=12070 1330 0 0 $X=11990 $Y=1080
X4 2 M3_M2_CDNS_1 $T=12670 2160 0 0 $X=12590 $Y=1910
X5 1 M2_M1_CDNS_2 $T=1170 1430 0 0 $X=1090 $Y=1180
X6 2 M2_M1_CDNS_2 $T=8020 1830 0 90 $X=7770 $Y=1750
X7 1 M2_M1_CDNS_2 $T=8650 1560 0 0 $X=8570 $Y=1310
X8 3 M2_M1_CDNS_2 $T=12070 1330 0 0 $X=11990 $Y=1080
X9 2 M2_M1_CDNS_2 $T=12670 2160 0 0 $X=12590 $Y=1910
X10 4 M4_M3_CDNS_3 $T=270 1810 0 180 $X=190 $Y=1560
X11 5 M4_M3_CDNS_3 $T=6460 1360 0 0 $X=6380 $Y=1110
X12 6 M4_M3_CDNS_3 $T=8070 1290 0 0 $X=7990 $Y=1040
X13 4 M4_M3_CDNS_3 $T=10010 1820 0 90 $X=9760 $Y=1740
X14 6 M4_M3_CDNS_3 $T=12110 1830 0 90 $X=11860 $Y=1750
X15 5 M4_M3_CDNS_3 $T=13590 1430 0 0 $X=13510 $Y=1180
X16 4 M2_M1_CDNS_4 $T=270 1810 0 180 $X=190 $Y=1560
X17 5 M2_M1_CDNS_4 $T=6460 1360 0 0 $X=6380 $Y=1110
X18 6 M2_M1_CDNS_4 $T=8070 1290 0 0 $X=7990 $Y=1040
X19 4 M2_M1_CDNS_4 $T=10010 1820 0 90 $X=9760 $Y=1740
X20 6 M2_M1_CDNS_4 $T=12110 1830 0 90 $X=11860 $Y=1750
X21 5 M2_M1_CDNS_4 $T=13590 1430 0 0 $X=13510 $Y=1180
X22 4 M3_M2_CDNS_5 $T=270 1810 0 180 $X=190 $Y=1560
X23 5 M3_M2_CDNS_5 $T=6460 1360 0 0 $X=6380 $Y=1110
X24 6 M3_M2_CDNS_5 $T=8070 1290 0 0 $X=7990 $Y=1040
X25 4 M3_M2_CDNS_5 $T=10010 1820 0 90 $X=9760 $Y=1740
X26 6 M3_M2_CDNS_5 $T=12110 1830 0 90 $X=11860 $Y=1750
X27 5 M3_M2_CDNS_5 $T=13590 1430 0 0 $X=13510 $Y=1180
X28 7 8 1 4 9 15 NAND2_1X $T=8400 -10 0 0 $X=8400 $Y=0
X29 7 8 9 6 3 16 NAND2_1X $T=10400 -10 0 0 $X=10400 $Y=0
X30 7 8 5 2 6 17 NAND2_2X $T=6400 0 0 0 $X=6400 $Y=0
X31 4 1 7 8 5 11 12 22 18 19 XOR2_1X $T=0 0 0 0 $X=0 $Y=0
X32 2 5 7 8 10 13 14 23 20 21 XOR2_1X $T=12400 0 0 0 $X=12400 $Y=0
M0 11 4 7 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=17.6861 scb=0.0184591 scc=0.000433664 $X=650 $Y=2490 $dt=1
M1 12 1 7 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.886 scb=0.00790338 scc=9.25552e-05 $X=1580 $Y=2490 $dt=1
M2 5 12 22 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=4880 $Y=2500 $dt=1
M3 7 4 22 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=5810 $Y=2500 $dt=1
M4 13 2 7 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=13050 $Y=2490 $dt=1
M5 14 5 7 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=13980 $Y=2490 $dt=1
M6 10 14 23 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6998 scb=0.00776618 scc=8.8963e-05 $X=17280 $Y=2500 $dt=1
M7 7 2 23 7 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.8514 scb=0.0153841 scc=0.000245782 $X=18210 $Y=2500 $dt=1
.ends 1_bit_Full_Adder_ver1
