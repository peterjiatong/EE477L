* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 10badder                                     *
* Netlisted  : Sun Nov 17 17:58:28 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_8                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_8 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_9                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_9 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_10                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_10 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_11                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_11 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_12                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_12 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_13                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_13 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_14                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_14 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_16                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_16 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_17                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_17 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_19                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_19 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_20                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_20 1 2 3
*.DEVICECLIMB
** N=3 EP=3 FDC=0
.ends nmos1v_CDNS_20

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_21                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_21 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_21

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_22                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_22 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_23                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_23 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_23

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_24                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_24 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_24

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=12
X0 7 M2_M1_CDNS_3 $T=250 -3000 0 0 $X=170 $Y=-3250
X1 7 M2_M1_CDNS_3 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X2 7 M1_PO_CDNS_8 $T=250 -3000 0 0 $X=150 $Y=-3250
X3 7 M1_PO_CDNS_8 $T=2620 -2730 0 0 $X=2520 $Y=-2980
X4 7 M3_M2_CDNS_9 $T=250 -3000 0 0 $X=170 $Y=-3250
X5 7 M3_M2_CDNS_9 $T=960 -2040 0 0 $X=880 $Y=-2290
X6 7 M3_M2_CDNS_9 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X7 1 M2_M1_CDNS_10 $T=1300 -3500 0 0 $X=1220 $Y=-3750
X8 1 M2_M1_CDNS_10 $T=2660 -4240 0 0 $X=2580 $Y=-4490
X9 1 M1_PO_CDNS_11 $T=1300 -3500 0 0 $X=1200 $Y=-3750
X10 1 M1_PO_CDNS_11 $T=2660 -4240 0 0 $X=2560 $Y=-4490
X11 7 M2_M1_CDNS_12 $T=960 -2040 0 0 $X=880 $Y=-2290
X12 1 M1_PO_CDNS_13 $T=680 -3550 0 0 $X=580 $Y=-3670
X13 4 M1_PO_CDNS_13 $T=1300 -2090 0 0 $X=1200 $Y=-2210
X14 5 M1_PO_CDNS_13 $T=4040 -3180 0 0 $X=3940 $Y=-3300
X15 8 M1_PO_CDNS_13 $T=4300 -3670 0 90 $X=4180 $Y=-3770
X16 3 8 6 2 3 pmos1v_CDNS_16 $T=4580 -3180 0 0 $X=4160 $Y=-3380
X17 2 6 8 2 nmos1v_CDNS_17 $T=4580 -4500 0 0 $X=4160 $Y=-4700
X18 3 1 7 2 3 pmos1v_CDNS_19 $T=750 -2850 0 0 $X=330 $Y=-3050
X19 2 7 1 nmos1v_CDNS_20 $T=750 -4370 0 0 $X=330 $Y=-4570
X20 2 7 9 2 nmos1v_CDNS_21 $T=1990 -4420 0 0 $X=1790 $Y=-4620
X21 8 5 10 2 nmos1v_CDNS_21 $T=3370 -4430 0 0 $X=3170 $Y=-4630
X22 8 4 9 2 nmos1v_CDNS_22 $T=1780 -4420 0 0 $X=1360 $Y=-4620
X23 2 1 10 2 nmos1v_CDNS_22 $T=3160 -4430 0 0 $X=2740 $Y=-4630
X24 3 1 11 2 3 pmos1v_CDNS_23 $T=1990 -3120 0 0 $X=1790 $Y=-3320
X25 8 5 12 2 3 pmos1v_CDNS_23 $T=3370 -3190 0 0 $X=3170 $Y=-3390
X26 8 4 11 2 3 pmos1v_CDNS_24 $T=1780 -3120 0 0 $X=1360 $Y=-3320
X27 3 7 12 2 3 pmos1v_CDNS_24 $T=3160 -3190 0 0 $X=2740 $Y=-3390
M0 7 1 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=750 $Y=-4370 $dt=0
M1 9 4 8 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1780 $Y=-4420 $dt=0
M2 2 7 9 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1990 $Y=-4420 $dt=0
M3 10 1 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3160 $Y=-4430 $dt=0
M4 8 5 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3370 $Y=-4430 $dt=0
M5 6 8 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=4580 $Y=-4500 $dt=0
M6 7 1 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=750 $Y=-2850 $dt=1
M7 11 4 8 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1780 $Y=-3120 $dt=1
M8 3 1 11 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1990 $Y=-3120 $dt=1
M9 12 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3160 $Y=-3190 $dt=1
M10 8 5 12 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3370 $Y=-3190 $dt=1
M11 6 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.2373 scb=0.0194294 scc=0.00149528 $X=4580 $Y=-3180 $dt=1
.ends MUX_2to1___2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_27                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_27 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_27

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_1X_small                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_27 $T=-310 120 0 0 $X=-430 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1000 $Y=830 $dt=0
M1 4 5 6 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1210 $Y=830 $dt=0
.ends NAND_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR1 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=6
X0 6 M2_M1_CDNS_5 $T=1210 1480 0 90 $X=1080 $Y=1400
X1 7 M2_M1_CDNS_5 $T=2250 1860 0 90 $X=2120 $Y=1780
X2 6 M2_M1_CDNS_5 $T=2950 1480 0 90 $X=2820 $Y=1400
X3 8 M2_M1_CDNS_5 $T=3370 650 0 0 $X=3290 $Y=520
X4 9 M2_M1_CDNS_5 $T=3370 3080 0 0 $X=3290 $Y=2950
X5 9 M2_M1_CDNS_5 $T=3930 3080 0 0 $X=3850 $Y=2950
X6 7 M2_M1_CDNS_5 $T=4680 1860 0 90 $X=4550 $Y=1780
X7 9 M2_M1_CDNS_5 $T=4890 3070 0 0 $X=4810 $Y=2940
X8 8 M2_M1_CDNS_5 $T=5840 640 0 0 $X=5760 $Y=510
X9 9 M2_M1_CDNS_5 $T=6260 3080 0 0 $X=6180 $Y=2950
X10 6 M1_PO_CDNS_13 $T=4020 1500 0 90 $X=3900 $Y=1400
X11 7 M1_PO_CDNS_13 $T=5020 1730 0 90 $X=4900 $Y=1630
X12 1 4 9 2 1 pmos1v_CDNS_16 $T=3120 2080 0 0 $X=2700 $Y=1880
X13 9 6 5 2 1 pmos1v_CDNS_16 $T=4090 2140 0 0 $X=3670 $Y=1940
X14 9 7 5 2 1 pmos1v_CDNS_16 $T=5050 2140 0 0 $X=4630 $Y=1940
X15 1 3 9 2 1 pmos1v_CDNS_16 $T=6010 2140 0 0 $X=5590 $Y=1940
X16 2 8 4 2 nmos1v_CDNS_17 $T=3120 780 0 0 $X=2700 $Y=580
X17 10 5 6 2 nmos1v_CDNS_17 $T=4090 760 0 0 $X=3670 $Y=560
X18 10 2 7 2 nmos1v_CDNS_17 $T=5050 770 0 0 $X=4630 $Y=570
X19 8 5 3 2 nmos1v_CDNS_17 $T=6010 770 0 0 $X=5590 $Y=570
X20 1 3 6 2 1 pmos1v_CDNS_19 $T=830 2320 0 0 $X=410 $Y=2120
X21 1 4 7 2 1 pmos1v_CDNS_19 $T=1790 2320 0 0 $X=1370 $Y=2120
X22 2 6 3 nmos1v_CDNS_20 $T=830 840 0 0 $X=410 $Y=640
X23 2 7 4 nmos1v_CDNS_20 $T=1790 840 0 0 $X=1370 $Y=640
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=830 $Y=840 $dt=0
M1 7 4 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1790 $Y=840 $dt=0
M2 8 4 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=3120 $Y=780 $dt=0
M3 5 6 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4126 scb=0.0095497 scc=0.000351079 $X=4090 $Y=760 $dt=0
M4 2 7 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=5050 $Y=770 $dt=0
M5 5 3 8 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=6010 $Y=770 $dt=0
.ends XOR1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_2X_small1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_2X_small1 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_27 $T=130 160 0 0 $X=10 $Y=20
M0 6 4 2 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=7.66878 scb=0.00580736 scc=7.77234e-05 $X=940 $Y=890 $dt=0
M1 3 5 6 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=11.676 scb=0.0124835 scc=0.000479408 $X=940 $Y=1100 $dt=0
.ends NAND_2X_small1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder1_small                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder1_small 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 22 23
*.DEVICECLIMB
** N=23 EP=16 FDC=18
X0 1 M2_M1_CDNS_3 $T=590 2080 0 90 $X=340 $Y=2000
X1 2 M2_M1_CDNS_3 $T=2300 3150 0 90 $X=2050 $Y=3070
X2 1 M2_M1_CDNS_3 $T=17380 1890 0 0 $X=17300 $Y=1640
X3 2 M2_M1_CDNS_3 $T=19040 3010 0 0 $X=18960 $Y=2760
X4 8 M2_M1_CDNS_5 $T=6580 1900 0 0 $X=6500 $Y=1770
X5 9 M2_M1_CDNS_5 $T=15190 1730 0 90 $X=15060 $Y=1650
X6 1 M1_PO_CDNS_8 $T=590 2080 0 90 $X=340 $Y=1980
X7 2 M1_PO_CDNS_8 $T=2300 3150 0 90 $X=2050 $Y=3050
X8 1 M1_PO_CDNS_8 $T=17380 1890 0 0 $X=17280 $Y=1640
X9 2 M1_PO_CDNS_8 $T=19040 3010 0 0 $X=18940 $Y=2760
X10 1 M3_M2_CDNS_9 $T=590 2080 0 90 $X=340 $Y=2000
X11 2 M3_M2_CDNS_9 $T=2300 3150 0 90 $X=2050 $Y=3070
X12 1 M3_M2_CDNS_9 $T=17380 1890 0 0 $X=17300 $Y=1640
X13 2 M3_M2_CDNS_9 $T=19040 3010 0 0 $X=18960 $Y=2760
X14 8 M2_M1_CDNS_10 $T=8510 1970 0 0 $X=8430 $Y=1720
X15 8 M2_M1_CDNS_10 $T=16110 1570 0 0 $X=16030 $Y=1320
X16 9 M2_M1_CDNS_10 $T=20260 1840 0 0 $X=20180 $Y=1590
X17 8 M1_PO_CDNS_11 $T=8510 1970 0 0 $X=8410 $Y=1720
X18 8 M1_PO_CDNS_11 $T=16110 1570 0 0 $X=16010 $Y=1320
X19 9 M1_PO_CDNS_11 $T=20260 1840 0 0 $X=20160 $Y=1590
X20 1 M1_PO_CDNS_13 $T=690 1610 0 0 $X=590 $Y=1490
X21 2 M1_PO_CDNS_13 $T=1650 1990 0 0 $X=1550 $Y=1870
X22 5 M1_PO_CDNS_13 $T=7590 1960 0 0 $X=7490 $Y=1840
X23 10 M1_PO_CDNS_13 $T=19320 1680 0 0 $X=19220 $Y=1560
X24 8 M3_M2_CDNS_14 $T=6970 950 0 0 $X=6890 $Y=820
X25 8 M3_M2_CDNS_14 $T=14100 570 0 90 $X=13970 $Y=490
X26 3 4 1 10 2 20 NAND_1X_small $T=16970 30 0 0 $X=16540 $Y=10
X27 3 4 9 7 10 21 NAND_1X_small $T=19810 30 0 0 $X=19380 $Y=10
X28 3 4 9 5 8 19 NAND_2X_small1 $T=13690 -10 0 0 $X=13700 $Y=10
X29 3 4 1 2 8 11 12 15 22 16 XOR1 $T=-40 30 0 0 $X=20 $Y=10
X30 3 4 5 8 6 13 14 17 23 18 XOR1 $T=6800 30 0 0 $X=6860 $Y=10
.ends full_adder1_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FA_4bit                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FA_4bit 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19
** N=83 EP=19 FDC=144
X0 17 M4_M3_CDNS_1 $T=14030 6120 0 0 $X=13950 $Y=5870
X1 18 M4_M3_CDNS_1 $T=16960 11880 0 0 $X=16880 $Y=11630
X2 17 M4_M3_CDNS_1 $T=19730 4760 0 0 $X=19650 $Y=4510
X3 18 M4_M3_CDNS_1 $T=22610 11350 0 0 $X=22530 $Y=11100
X4 17 M3_M2_CDNS_2 $T=14030 6120 0 0 $X=13950 $Y=5870
X5 18 M3_M2_CDNS_2 $T=16960 11880 0 0 $X=16880 $Y=11630
X6 18 M3_M2_CDNS_2 $T=22610 11350 0 0 $X=22530 $Y=11100
X7 17 M2_M1_CDNS_3 $T=14030 6120 0 0 $X=13950 $Y=5870
X8 18 M2_M1_CDNS_3 $T=16960 11880 0 0 $X=16880 $Y=11630
X9 19 M2_M1_CDNS_3 $T=18840 8310 0 0 $X=18760 $Y=8060
X10 18 M2_M1_CDNS_3 $T=22610 11350 0 0 $X=22530 $Y=11100
X11 1 M2_M1_CDNS_5 $T=-80 3540 0 0 $X=-160 $Y=3410
X12 1 M2_M1_CDNS_5 $T=-80 10890 0 0 $X=-160 $Y=10760
X13 17 M2_M1_CDNS_5 $T=21770 2020 0 0 $X=21690 $Y=1890
X14 19 M2_M1_CDNS_5 $T=21770 5100 0 0 $X=21690 $Y=4970
X15 17 M1_PO_CDNS_8 $T=14030 6120 0 0 $X=13930 $Y=5870
X16 18 M1_PO_CDNS_8 $T=16960 11880 0 0 $X=16860 $Y=11630
X17 19 M1_PO_CDNS_8 $T=18840 8310 0 0 $X=18740 $Y=8060
X18 19 M3_M2_CDNS_9 $T=18840 8310 0 0 $X=18760 $Y=8060
X19 19 M3_M2_CDNS_14 $T=21980 9220 0 0 $X=21900 $Y=9090
X20 3 2 1 10 11 12 17 43 46 47
+ 41 42 44 45 82 83 full_adder1_small $T=-90 -130 0 0 $X=-70 $Y=-120
X21 5 4 1 10 17 13 19 36 39 40
+ 34 35 37 38 80 81 full_adder1_small $T=-90 7250 1 0 $X=-70 $Y=3440
X22 7 6 1 10 19 14 18 29 32 33
+ 27 28 30 31 78 79 full_adder1_small $T=-90 7190 0 0 $X=-70 $Y=7200
X23 9 8 1 10 18 15 16 22 25 26
+ 20 21 23 24 76 77 full_adder1_small $T=-90 14570 1 0 $X=-70 $Y=10760
M0 41 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=2220 $dt=1
M1 34 5 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=4420 $dt=1
M2 27 7 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=9540 $dt=1
M3 20 9 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=11740 $dt=1
M4 42 2 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=2220 $dt=1
M5 35 4 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=4420 $dt=1
M6 28 6 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=9540 $dt=1
M7 21 8 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=11740 $dt=1
M8 82 2 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=1980 $dt=1
M9 80 4 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=4180 $dt=1
M10 78 6 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=9300 $dt=1
M11 76 8 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=11500 $dt=1
M12 43 41 82 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=2040 $dt=1
M13 36 34 80 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=4120 $dt=1
M14 29 27 78 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=9360 $dt=1
M15 22 20 76 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=11440 $dt=1
M16 43 42 82 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=2040 $dt=1
M17 36 35 80 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=4120 $dt=1
M18 29 28 78 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=9360 $dt=1
M19 22 21 76 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=11440 $dt=1
M20 82 3 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=2040 $dt=1
M21 80 5 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=4120 $dt=1
M22 78 7 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=9360 $dt=1
M23 76 9 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=11440 $dt=1
M24 44 11 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=2220 $dt=1
M25 37 17 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=4420 $dt=1
M26 30 19 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=9540 $dt=1
M27 23 18 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=11740 $dt=1
M28 45 43 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=2220 $dt=1
M29 38 36 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=4420 $dt=1
M30 31 29 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=9540 $dt=1
M31 24 22 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=11740 $dt=1
M32 83 43 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=1980 $dt=1
M33 81 36 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=4180 $dt=1
M34 79 29 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=9300 $dt=1
M35 77 22 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=11500 $dt=1
M36 12 44 83 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=2040 $dt=1
M37 13 37 81 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=4120 $dt=1
M38 14 30 79 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=9360 $dt=1
M39 15 23 77 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=11440 $dt=1
M40 12 45 83 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=2040 $dt=1
M41 13 38 81 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=4120 $dt=1
M42 14 31 79 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=9360 $dt=1
M43 15 24 77 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=11440 $dt=1
M44 83 11 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=2040 $dt=1
M45 81 17 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=4120 $dt=1
M46 79 19 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=9360 $dt=1
M47 77 18 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=11440 $dt=1
M48 46 11 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=2010 $dt=1
M49 39 17 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=4150 $dt=1
M50 32 19 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=9330 $dt=1
M51 25 18 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=11470 $dt=1
M52 1 43 46 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=2010 $dt=1
M53 1 36 39 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=4150 $dt=1
M54 1 29 32 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=9330 $dt=1
M55 1 22 25 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=11470 $dt=1
M56 47 3 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=2230 $dt=1
M57 40 5 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=4410 $dt=1
M58 33 7 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=9550 $dt=1
M59 26 9 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=11730 $dt=1
M60 1 2 47 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=2230 $dt=1
M61 1 4 40 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=4410 $dt=1
M62 1 6 33 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=9550 $dt=1
M63 1 8 26 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=11730 $dt=1
M64 17 46 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=2230 $dt=1
M65 19 39 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=4410 $dt=1
M66 18 32 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=9550 $dt=1
M67 16 25 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=11730 $dt=1
M68 1 47 17 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=2230 $dt=1
M69 1 40 19 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=4410 $dt=1
M70 1 33 18 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=9550 $dt=1
M71 1 26 16 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=11730 $dt=1
.ends FA_4bit

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small 1 2 3 4
** N=4 EP=4 FDC=2
X0 1 M1_PO_CDNS_13 $T=950 1780 0 90 $X=830 $Y=1680
X1 2 1 4 3 2 pmos1v_CDNS_19 $T=1070 2220 0 0 $X=650 $Y=2020
X2 3 4 1 nmos1v_CDNS_20 $T=1070 980 0 0 $X=650 $Y=780
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7353 scb=0.0117274 scc=0.000445561 $X=1070 $Y=980 $dt=0
M1 4 1 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8675 scb=0.0146094 scc=0.000688105 $X=1070 $Y=2220 $dt=1
.ends INV_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 10badder                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 10badder 6 51 52 53 54 55 56 57 58 59
+ 47 50 38 21 39 40 41 23 42 43
+ 44 46 48 30 17 22 18 31 19 24
+ 20 45 49 25
** N=267 EP=34 FDC=516
X0 1 M4_M3_CDNS_1 $T=51080 34160 0 0 $X=51000 $Y=33910
X1 2 M4_M3_CDNS_1 $T=56340 32800 0 0 $X=56260 $Y=32550
X2 3 M4_M3_CDNS_1 $T=56340 47440 0 0 $X=56260 $Y=47190
X3 4 M4_M3_CDNS_1 $T=57240 50840 0 0 $X=57160 $Y=50590
X4 5 M4_M3_CDNS_1 $T=72650 52420 0 90 $X=72400 $Y=52340
X5 1 M4_M3_CDNS_1 $T=78550 36430 0 0 $X=78470 $Y=36180
X6 5 M4_M3_CDNS_1 $T=79400 52420 0 90 $X=79150 $Y=52340
X7 2 M4_M3_CDNS_1 $T=86760 34460 0 0 $X=86680 $Y=34210
X8 3 M4_M3_CDNS_1 $T=86760 49100 0 0 $X=86680 $Y=48850
X9 1 M3_M2_CDNS_2 $T=51080 34160 0 0 $X=51000 $Y=33910
X10 2 M3_M2_CDNS_2 $T=56340 32800 0 0 $X=56260 $Y=32550
X11 3 M3_M2_CDNS_2 $T=56340 47440 0 0 $X=56260 $Y=47190
X12 4 M3_M2_CDNS_2 $T=57240 50840 0 0 $X=57160 $Y=50590
X13 5 M3_M2_CDNS_2 $T=72650 52420 0 90 $X=72400 $Y=52340
X14 1 M3_M2_CDNS_2 $T=78550 36430 0 0 $X=78470 $Y=36180
X15 5 M3_M2_CDNS_2 $T=79400 52420 0 90 $X=79150 $Y=52340
X16 2 M3_M2_CDNS_2 $T=86760 34460 0 0 $X=86680 $Y=34210
X17 3 M3_M2_CDNS_2 $T=86760 49100 0 0 $X=86680 $Y=48850
X18 1 M2_M1_CDNS_3 $T=51080 34160 0 0 $X=51000 $Y=33910
X19 6 M2_M1_CDNS_3 $T=52330 32180 0 90 $X=52080 $Y=32100
X20 1 M2_M1_CDNS_3 $T=52330 46820 0 90 $X=52080 $Y=46740
X21 7 M2_M1_CDNS_3 $T=54270 29810 0 90 $X=54020 $Y=29730
X22 8 M2_M1_CDNS_3 $T=54270 44450 0 90 $X=54020 $Y=44370
X23 9 M2_M1_CDNS_3 $T=55540 26280 0 0 $X=55460 $Y=26030
X24 10 M2_M1_CDNS_3 $T=55540 40920 0 0 $X=55460 $Y=40670
X25 11 M2_M1_CDNS_3 $T=55730 21200 0 90 $X=55480 $Y=21120
X26 12 M2_M1_CDNS_3 $T=55730 35840 0 90 $X=55480 $Y=35760
X27 13 M2_M1_CDNS_3 $T=56210 23810 0 90 $X=55960 $Y=23730
X28 14 M2_M1_CDNS_3 $T=56210 38450 0 90 $X=55960 $Y=38370
X29 15 M2_M1_CDNS_3 $T=56050 31070 0 0 $X=55970 $Y=30820
X30 16 M2_M1_CDNS_3 $T=56050 45710 0 0 $X=55970 $Y=45460
X31 2 M2_M1_CDNS_3 $T=56340 32800 0 0 $X=56260 $Y=32550
X32 3 M2_M1_CDNS_3 $T=56340 47440 0 0 $X=56260 $Y=47190
X33 4 M2_M1_CDNS_3 $T=57240 50840 0 0 $X=57160 $Y=50590
X34 17 M2_M1_CDNS_3 $T=57660 26200 0 90 $X=57410 $Y=26120
X35 18 M2_M1_CDNS_3 $T=57660 33520 0 90 $X=57410 $Y=33440
X36 19 M2_M1_CDNS_3 $T=57660 40840 0 90 $X=57410 $Y=40760
X37 20 M2_M1_CDNS_3 $T=57660 48160 0 90 $X=57410 $Y=48080
X38 21 M2_M1_CDNS_3 $T=57670 22770 0 90 $X=57420 $Y=22690
X39 22 M2_M1_CDNS_3 $T=57670 30070 0 90 $X=57420 $Y=29990
X40 23 M2_M1_CDNS_3 $T=57670 37410 0 90 $X=57420 $Y=37330
X41 24 M2_M1_CDNS_3 $T=57670 44710 0 90 $X=57420 $Y=44630
X42 5 M2_M1_CDNS_3 $T=72650 52420 0 90 $X=72400 $Y=52340
X43 1 M2_M1_CDNS_3 $T=78550 36430 0 0 $X=78470 $Y=36180
X44 5 M2_M1_CDNS_3 $T=79400 52420 0 90 $X=79150 $Y=52340
X45 2 M2_M1_CDNS_3 $T=86760 34460 0 0 $X=86680 $Y=34210
X46 3 M2_M1_CDNS_3 $T=86760 49100 0 0 $X=86680 $Y=48850
X47 25 M2_M1_CDNS_5 $T=50480 50560 0 0 $X=50400 $Y=50430
X48 25 M2_M1_CDNS_5 $T=51590 45750 0 90 $X=51460 $Y=45670
X49 26 M2_M1_CDNS_5 $T=53210 27000 0 0 $X=53130 $Y=26870
X50 27 M2_M1_CDNS_5 $T=53210 41640 0 0 $X=53130 $Y=41510
X51 28 M2_M1_CDNS_5 $T=53230 23140 0 0 $X=53150 $Y=23010
X52 29 M2_M1_CDNS_5 $T=53230 37780 0 0 $X=53150 $Y=37650
X53 25 M2_M1_CDNS_5 $T=62920 24380 0 0 $X=62840 $Y=24250
X54 25 M2_M1_CDNS_5 $T=62920 39020 0 0 $X=62840 $Y=38890
X55 25 M2_M1_CDNS_5 $T=62930 31710 0 0 $X=62850 $Y=31580
X56 25 M2_M1_CDNS_5 $T=62930 46350 0 0 $X=62850 $Y=46220
X57 6 M1_PO_CDNS_8 $T=52330 32180 0 90 $X=52080 $Y=32080
X58 1 M1_PO_CDNS_8 $T=52330 46820 0 90 $X=52080 $Y=46720
X59 7 M1_PO_CDNS_8 $T=54270 29810 0 90 $X=54020 $Y=29710
X60 8 M1_PO_CDNS_8 $T=54270 44450 0 90 $X=54020 $Y=44350
X61 9 M1_PO_CDNS_8 $T=55540 26280 0 0 $X=55440 $Y=26030
X62 10 M1_PO_CDNS_8 $T=55540 40920 0 0 $X=55440 $Y=40670
X63 11 M1_PO_CDNS_8 $T=55730 21200 0 90 $X=55480 $Y=21100
X64 12 M1_PO_CDNS_8 $T=55730 35840 0 90 $X=55480 $Y=35740
X65 15 M1_PO_CDNS_8 $T=56050 31070 0 0 $X=55950 $Y=30820
X66 16 M1_PO_CDNS_8 $T=56050 45710 0 0 $X=55950 $Y=45460
X67 13 M1_PO_CDNS_8 $T=56210 23810 0 90 $X=55960 $Y=23710
X68 14 M1_PO_CDNS_8 $T=56210 38450 0 90 $X=55960 $Y=38350
X69 2 M1_PO_CDNS_8 $T=56340 32800 0 0 $X=56240 $Y=32550
X70 3 M1_PO_CDNS_8 $T=56340 47440 0 0 $X=56240 $Y=47190
X71 17 M1_PO_CDNS_8 $T=57660 26200 0 90 $X=57410 $Y=26100
X72 18 M1_PO_CDNS_8 $T=57660 33520 0 90 $X=57410 $Y=33420
X73 19 M1_PO_CDNS_8 $T=57660 40840 0 90 $X=57410 $Y=40740
X74 20 M1_PO_CDNS_8 $T=57660 48160 0 90 $X=57410 $Y=48060
X75 21 M1_PO_CDNS_8 $T=57670 22770 0 90 $X=57420 $Y=22670
X76 22 M1_PO_CDNS_8 $T=57670 30070 0 90 $X=57420 $Y=29970
X77 23 M1_PO_CDNS_8 $T=57670 37410 0 90 $X=57420 $Y=37310
X78 24 M1_PO_CDNS_8 $T=57670 44710 0 90 $X=57420 $Y=44610
X79 1 M1_PO_CDNS_8 $T=78550 36430 0 0 $X=78450 $Y=36180
X80 6 M3_M2_CDNS_9 $T=52330 32180 0 90 $X=52080 $Y=32100
X81 1 M3_M2_CDNS_9 $T=52330 46820 0 90 $X=52080 $Y=46740
X82 9 M3_M2_CDNS_9 $T=53480 29020 0 0 $X=53400 $Y=28770
X83 10 M3_M2_CDNS_9 $T=53480 43660 0 0 $X=53400 $Y=43410
X84 7 M3_M2_CDNS_9 $T=54270 29810 0 90 $X=54020 $Y=29730
X85 8 M3_M2_CDNS_9 $T=54270 44450 0 90 $X=54020 $Y=44370
X86 9 M3_M2_CDNS_9 $T=55540 26280 0 0 $X=55460 $Y=26030
X87 10 M3_M2_CDNS_9 $T=55540 40920 0 0 $X=55460 $Y=40670
X88 11 M3_M2_CDNS_9 $T=55730 21200 0 90 $X=55480 $Y=21120
X89 12 M3_M2_CDNS_9 $T=55730 35840 0 90 $X=55480 $Y=35760
X90 13 M3_M2_CDNS_9 $T=56210 23810 0 90 $X=55960 $Y=23730
X91 14 M3_M2_CDNS_9 $T=56210 38450 0 90 $X=55960 $Y=38370
X92 15 M3_M2_CDNS_9 $T=56050 31070 0 0 $X=55970 $Y=30820
X93 16 M3_M2_CDNS_9 $T=56050 45710 0 0 $X=55970 $Y=45460
X94 26 M3_M2_CDNS_9 $T=56240 34220 0 0 $X=56160 $Y=33970
X95 27 M3_M2_CDNS_9 $T=56240 48860 0 0 $X=56160 $Y=48610
X96 17 M3_M2_CDNS_9 $T=57660 26200 0 90 $X=57410 $Y=26120
X97 18 M3_M2_CDNS_9 $T=57660 33520 0 90 $X=57410 $Y=33440
X98 19 M3_M2_CDNS_9 $T=57660 40840 0 90 $X=57410 $Y=40760
X99 20 M3_M2_CDNS_9 $T=57660 48160 0 90 $X=57410 $Y=48080
X100 21 M3_M2_CDNS_9 $T=57670 22770 0 90 $X=57420 $Y=22690
X101 22 M3_M2_CDNS_9 $T=57670 30070 0 90 $X=57420 $Y=29990
X102 23 M3_M2_CDNS_9 $T=57670 37410 0 90 $X=57420 $Y=37330
X103 24 M3_M2_CDNS_9 $T=57670 44710 0 90 $X=57420 $Y=44630
X104 15 M3_M2_CDNS_9 $T=62950 31240 0 90 $X=62700 $Y=31160
X105 16 M3_M2_CDNS_9 $T=62950 45880 0 90 $X=62700 $Y=45800
X106 13 M3_M2_CDNS_9 $T=63400 23460 0 0 $X=63320 $Y=23210
X107 14 M3_M2_CDNS_9 $T=63400 38100 0 0 $X=63320 $Y=37850
X108 11 M3_M2_CDNS_9 $T=63720 21760 0 0 $X=63640 $Y=21510
X109 12 M3_M2_CDNS_9 $T=63720 36400 0 0 $X=63640 $Y=36150
X110 7 M3_M2_CDNS_9 $T=63820 29420 0 0 $X=63740 $Y=29170
X111 8 M3_M2_CDNS_9 $T=63820 44060 0 0 $X=63740 $Y=43810
X112 28 M2_M1_CDNS_10 $T=53520 24980 0 90 $X=53270 $Y=24900
X113 29 M2_M1_CDNS_10 $T=53520 39620 0 90 $X=53270 $Y=39540
X114 30 M2_M1_CDNS_10 $T=64110 23330 0 0 $X=64030 $Y=23080
X115 31 M2_M1_CDNS_10 $T=64110 37970 0 0 $X=64030 $Y=37720
X116 30 M2_M1_CDNS_10 $T=65950 23850 0 90 $X=65700 $Y=23770
X117 31 M2_M1_CDNS_10 $T=65950 38490 0 90 $X=65700 $Y=38410
X118 6 M2_M1_CDNS_10 $T=78510 22370 0 0 $X=78430 $Y=22120
X119 28 M1_PO_CDNS_11 $T=53520 24980 0 90 $X=53270 $Y=24880
X120 29 M1_PO_CDNS_11 $T=53520 39620 0 90 $X=53270 $Y=39520
X121 30 M1_PO_CDNS_11 $T=64110 23330 0 0 $X=64010 $Y=23080
X122 31 M1_PO_CDNS_11 $T=64110 37970 0 0 $X=64010 $Y=37720
X123 30 M1_PO_CDNS_11 $T=65950 23850 0 90 $X=65700 $Y=23750
X124 31 M1_PO_CDNS_11 $T=65950 38490 0 90 $X=65700 $Y=38390
X125 6 M1_PO_CDNS_11 $T=78510 22370 0 0 $X=78410 $Y=22120
X126 9 M2_M1_CDNS_12 $T=53480 29020 0 0 $X=53400 $Y=28770
X127 10 M2_M1_CDNS_12 $T=53480 43660 0 0 $X=53400 $Y=43410
X128 26 M2_M1_CDNS_12 $T=56240 34220 0 0 $X=56160 $Y=33970
X129 27 M2_M1_CDNS_12 $T=56240 48860 0 0 $X=56160 $Y=48610
X130 15 M2_M1_CDNS_12 $T=62950 31240 0 90 $X=62700 $Y=31160
X131 16 M2_M1_CDNS_12 $T=62950 45880 0 90 $X=62700 $Y=45800
X132 13 M2_M1_CDNS_12 $T=63400 23460 0 0 $X=63320 $Y=23210
X133 14 M2_M1_CDNS_12 $T=63400 38100 0 0 $X=63320 $Y=37850
X134 11 M2_M1_CDNS_12 $T=63720 21760 0 0 $X=63640 $Y=21510
X135 12 M2_M1_CDNS_12 $T=63720 36400 0 0 $X=63640 $Y=36150
X136 7 M2_M1_CDNS_12 $T=63820 29420 0 0 $X=63740 $Y=29170
X137 8 M2_M1_CDNS_12 $T=63820 44060 0 0 $X=63740 $Y=43810
X138 32 M1_PO_CDNS_13 $T=53270 31100 0 0 $X=53170 $Y=30980
X139 33 M1_PO_CDNS_13 $T=53270 45740 0 0 $X=53170 $Y=45620
X140 34 M1_PO_CDNS_13 $T=53550 23450 0 0 $X=53450 $Y=23330
X141 35 M1_PO_CDNS_13 $T=53550 38090 0 0 $X=53450 $Y=37970
X142 36 M1_PO_CDNS_13 $T=53840 25910 0 0 $X=53740 $Y=25790
X143 37 M1_PO_CDNS_13 $T=53840 40550 0 0 $X=53740 $Y=40430
X144 26 M3_M2_CDNS_14 $T=50730 34460 0 0 $X=50650 $Y=34330
X145 27 M3_M2_CDNS_14 $T=50800 49100 0 0 $X=50720 $Y=48970
X146 6 M3_M2_CDNS_14 $T=51610 22610 0 0 $X=51530 $Y=22480
X147 26 38 25 2 6 1 60 61 156 157
+ 252 253 MUX_2to1___2X $T=56190 30160 0 180 $X=50640 $Y=31580
X148 27 38 25 3 1 4 62 63 158 159
+ 254 255 MUX_2to1___2X $T=56190 44800 0 180 $X=50640 $Y=46220
X149 25 38 11 34 13 160 NAND_1X_small $T=53960 20720 0 0 $X=53530 $Y=20700
X150 25 38 9 36 28 161 NAND_1X_small $T=55940 28040 0 180 $X=53530 $Y=24260
X151 25 38 7 32 15 162 NAND_1X_small $T=53960 28040 0 0 $X=53530 $Y=28020
X152 25 38 12 35 14 163 NAND_1X_small $T=53960 35360 0 0 $X=53530 $Y=35340
X153 25 38 10 37 29 164 NAND_1X_small $T=55940 42680 0 180 $X=53530 $Y=38900
X154 25 38 8 33 16 165 NAND_1X_small $T=53960 42680 0 0 $X=53530 $Y=42660
X155 25 38 30 21 13 64 65 166 256 167 XOR1 $T=56070 20720 0 0 $X=56130 $Y=20700
X156 25 38 39 17 11 66 67 168 257 169 XOR1 $T=56070 28040 1 0 $X=56130 $Y=24260
X157 25 38 40 22 15 68 69 170 258 171 XOR1 $T=56070 28040 0 0 $X=56130 $Y=28020
X158 25 38 41 18 7 70 71 172 259 173 XOR1 $T=56070 35360 1 0 $X=56130 $Y=31580
X159 25 38 31 23 14 72 73 174 260 175 XOR1 $T=56070 35360 0 0 $X=56130 $Y=35340
X160 25 38 42 19 12 74 75 176 261 177 XOR1 $T=56070 42680 1 0 $X=56130 $Y=38900
X161 25 38 43 24 16 76 77 178 262 179 XOR1 $T=56070 42680 0 0 $X=56130 $Y=42660
X162 25 38 44 20 8 78 79 180 263 181 XOR1 $T=56070 50000 1 0 $X=56130 $Y=46220
X163 45 46 25 38 4 47 5 82 85 86
+ 80 81 83 84 264 265 full_adder1_small $T=50650 49970 0 0 $X=50670 $Y=49980
X164 48 49 25 38 5 50 51 89 92 93
+ 87 88 90 91 266 267 full_adder1_small $T=72610 49970 0 0 $X=72630 $Y=49980
X165 25 30 21 17 39 22 40 18 41 38
+ 6 52 53 54 55 2 114 115 116 FA_4bit $T=64900 20820 0 0 $X=64250 $Y=20700
X166 25 31 23 19 42 24 43 20 44 38
+ 1 56 57 58 59 3 145 146 147 FA_4bit $T=64900 35460 0 0 $X=64250 $Y=35340
X167 34 25 38 28 INV_1X_small $T=51530 20700 0 0 $X=51530 $Y=20700
X168 36 25 38 26 INV_1X_small $T=51530 28060 1 0 $X=51530 $Y=24260
X169 32 25 38 9 INV_1X_small $T=51530 28020 0 0 $X=51530 $Y=28020
X170 35 25 38 29 INV_1X_small $T=51530 35340 0 0 $X=51530 $Y=35340
X171 37 25 38 27 INV_1X_small $T=51530 42700 1 0 $X=51530 $Y=38900
X172 33 25 38 10 INV_1X_small $T=51530 42660 0 0 $X=51530 $Y=42660
M0 80 45 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6612 scb=0.0167915 scc=0.000377457 $X=51440 $Y=52320 $dt=1
M1 81 46 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.8911 scb=0.00996238 scc=0.000256798 $X=52400 $Y=52320 $dt=1
M2 264 46 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=53730 $Y=52080 $dt=1
M3 36 28 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=25230 $dt=1
M4 37 29 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=39870 $dt=1
M5 82 80 264 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=54700 $Y=52140 $dt=1
M6 34 11 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=23050 $dt=1
M7 32 7 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=30370 $dt=1
M8 35 12 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=37690 $dt=1
M9 33 8 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=45010 $dt=1
M10 25 9 36 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=25230 $dt=1
M11 25 10 37 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=39870 $dt=1
M12 25 13 34 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=23050 $dt=1
M13 25 15 32 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=30370 $dt=1
M14 25 14 35 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=37690 $dt=1
M15 25 16 33 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=45010 $dt=1
M16 82 81 264 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=55660 $Y=52140 $dt=1
M17 264 45 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=56620 $Y=52140 $dt=1
M18 64 30 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=23040 $dt=1
M19 66 39 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=25240 $dt=1
M20 68 40 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=30360 $dt=1
M21 70 41 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=32560 $dt=1
M22 72 31 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=37680 $dt=1
M23 74 42 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=39880 $dt=1
M24 76 43 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=45000 $dt=1
M25 78 44 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=47200 $dt=1
M26 65 21 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=23040 $dt=1
M27 67 17 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=25240 $dt=1
M28 69 22 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=30360 $dt=1
M29 71 18 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=32560 $dt=1
M30 73 23 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=37680 $dt=1
M31 75 19 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=39880 $dt=1
M32 77 24 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=45000 $dt=1
M33 79 20 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=47200 $dt=1
M34 83 4 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=58280 $Y=52320 $dt=1
M35 256 21 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=22800 $dt=1
M36 257 17 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=25000 $dt=1
M37 258 22 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=30120 $dt=1
M38 259 18 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=32320 $dt=1
M39 260 23 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=37440 $dt=1
M40 261 19 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=39640 $dt=1
M41 262 24 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=44760 $dt=1
M42 263 20 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=46960 $dt=1
M43 84 82 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=59240 $Y=52320 $dt=1
M44 13 64 256 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=22860 $dt=1
M45 11 66 257 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=24940 $dt=1
M46 15 68 258 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=30180 $dt=1
M47 7 70 259 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=32260 $dt=1
M48 14 72 260 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=37500 $dt=1
M49 12 74 261 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=39580 $dt=1
M50 16 76 262 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=44820 $dt=1
M51 8 78 263 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=46900 $dt=1
M52 265 82 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60570 $Y=52080 $dt=1
M53 13 65 256 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=22860 $dt=1
M54 11 67 257 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=24940 $dt=1
M55 15 69 258 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=30180 $dt=1
M56 7 71 259 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=32260 $dt=1
M57 14 73 260 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=37500 $dt=1
M58 12 75 261 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=39580 $dt=1
M59 16 77 262 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=44820 $dt=1
M60 8 79 263 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=46900 $dt=1
M61 47 83 265 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=61540 $Y=52140 $dt=1
M62 256 30 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=22860 $dt=1
M63 257 39 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=24940 $dt=1
M64 258 40 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=30180 $dt=1
M65 259 41 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=32260 $dt=1
M66 260 31 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=37500 $dt=1
M67 261 42 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=39580 $dt=1
M68 262 43 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=44820 $dt=1
M69 263 44 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=46900 $dt=1
M70 47 84 265 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=62500 $Y=52140 $dt=1
M71 265 4 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=63460 $Y=52140 $dt=1
M72 85 4 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65530 $Y=52110 $dt=1
M73 25 82 85 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65940 $Y=52110 $dt=1
M74 86 45 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68510 $Y=52330 $dt=1
M75 25 46 86 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68920 $Y=52330 $dt=1
M76 5 85 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71350 $Y=52330 $dt=1
M77 25 86 5 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71760 $Y=52330 $dt=1
M78 87 48 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=73400 $Y=52320 $dt=1
M79 88 49 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=74360 $Y=52320 $dt=1
M80 266 49 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=75690 $Y=52080 $dt=1
M81 89 87 266 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=76660 $Y=52140 $dt=1
M82 89 88 266 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=77620 $Y=52140 $dt=1
M83 266 48 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=78580 $Y=52140 $dt=1
M84 90 5 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=80240 $Y=52320 $dt=1
M85 91 89 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=81200 $Y=52320 $dt=1
M86 267 89 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=82530 $Y=52080 $dt=1
M87 50 90 267 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=83500 $Y=52140 $dt=1
M88 50 91 267 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=84460 $Y=52140 $dt=1
M89 267 5 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=85420 $Y=52140 $dt=1
M90 92 5 25 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87490 $Y=52110 $dt=1
M91 25 89 92 25 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87900 $Y=52110 $dt=1
M92 93 48 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90470 $Y=52330 $dt=1
M93 25 49 93 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90880 $Y=52330 $dt=1
M94 51 92 25 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=93310 $Y=52330 $dt=1
M95 25 93 51 25 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=93720 $Y=52330 $dt=1
.ends 10badder
