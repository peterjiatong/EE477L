* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : AND4_1x                                      *
* Netlisted  : Sun Nov  3 06:41:16 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_6                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_6 D_drain_1 2 3 4
** N=4 EP=4 FDC=1
M0 D_drain_1 2 3 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_7                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_7 S_source_0 2 3
** N=3 EP=3 FDC=1
M0 3 2 S_source_0 S_source_0 g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X in_b in_a out vdd! gnd!
*.DEVICECLIMB
** N=6 EP=5 FDC=2
X4 out in_b 6 gnd! nmos1v_CDNS_6 $T=830 720 0 0 $X=630 $Y=520
X5 gnd! in_a 6 nmos1v_CDNS_7 $T=620 720 0 0 $X=200 $Y=520
.ends NAND2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_8                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_8 S_source_0 D_drain_1 3
** N=3 EP=3 FDC=1
M0 D_drain_1 3 S_source_0 S_source_0 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6908 scb=0.0179614 scc=0.00130074 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X out in vdd! gnd!
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X1 gnd! out in nmos1v_CDNS_8 $T=1090 1110 0 0 $X=670 $Y=910
.ends INV_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND4_1x                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND4_1x A B C D OUT gnd! vdd!
** N=15 EP=7 FDC=18
X2 B A 4 vdd! gnd! NAND2_1X $T=0 -10 0 0 $X=0 $Y=0
X3 D C 9 vdd! gnd! NAND2_1X $T=4000 -10 0 0 $X=4000 $Y=0
X4 1 10 11 vdd! gnd! NAND2_1X $T=8000 -10 0 0 $X=8000 $Y=0
X5 1 4 vdd! gnd! INV_1X $T=1990 0 0 0 $X=2000 $Y=0
X6 10 9 vdd! gnd! INV_1X $T=5990 0 0 0 $X=6000 $Y=0
X7 OUT 11 vdd! gnd! INV_1X $T=9990 0 0 0 $X=10000 $Y=0
M0 4 A vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=29.8065 scb=0.0321965 scc=0.00263528 $X=620 $Y=2070 $dt=1
M1 vdd! B 4 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=24.1872 scb=0.0226978 scc=0.00220665 $X=1030 $Y=2070 $dt=1
M2 1 4 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=18.2452 scb=0.0177397 scc=0.00150411 $X=3080 $Y=2120 $dt=1
M3 9 C vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=4620 $Y=2070 $dt=1
M4 vdd! D 9 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=5030 $Y=2070 $dt=1
M5 10 9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=18.2452 scb=0.0177397 scc=0.00150411 $X=7080 $Y=2120 $dt=1
M6 11 10 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=8620 $Y=2070 $dt=1
M7 vdd! 1 11 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=9030 $Y=2070 $dt=1
M8 OUT 11 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=20.511 scb=0.0198276 scc=0.00151235 $X=11080 $Y=2120 $dt=1
.ends AND4_1x
