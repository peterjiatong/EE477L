* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : MUX_2to1___2X_forph2p2                       *
* Netlisted  : Sun Nov 24 15:20:42 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_8                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_8 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_9                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_9 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_11                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_11 1 2 3 4 5
** N=5 EP=5 FDC=1
M0 2 3 1 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.4542 scb=0.0129422 scc=0.000231427 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_12                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_12 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_13                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_13 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_14                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_14 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_15                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_15 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_16                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_16 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X_forph2p2                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X_forph2p2 2 3 1 8 7 6
** N=12 EP=6 FDC=12
X0 1 M2_M1_CDNS_1 $T=1480 1720 0 0 $X=1400 $Y=1470
X1 1 M2_M1_CDNS_1 $T=2840 980 0 0 $X=2760 $Y=730
X2 1 M1_PO_CDNS_2 $T=1480 1720 0 0 $X=1380 $Y=1470
X3 1 M1_PO_CDNS_2 $T=2840 980 0 0 $X=2740 $Y=730
X4 1 M1_PO_CDNS_3 $T=860 1670 0 0 $X=760 $Y=1550
X5 2 M1_PO_CDNS_3 $T=1480 3130 0 0 $X=1380 $Y=3010
X6 3 M1_PO_CDNS_3 $T=4220 2040 0 0 $X=4120 $Y=1920
X7 4 M1_PO_CDNS_3 $T=4480 1550 0 90 $X=4360 $Y=1450
X8 5 M3_M2_CDNS_5 $T=430 2220 0 0 $X=350 $Y=1970
X9 5 M3_M2_CDNS_5 $T=1140 3180 0 0 $X=1060 $Y=2930
X10 5 M3_M2_CDNS_5 $T=2800 2490 0 0 $X=2720 $Y=2240
X11 5 M2_M1_CDNS_6 $T=430 2220 0 0 $X=350 $Y=1970
X12 5 M2_M1_CDNS_6 $T=2800 2490 0 0 $X=2720 $Y=2240
X13 5 M1_PO_CDNS_7 $T=430 2220 0 0 $X=330 $Y=1970
X14 5 M1_PO_CDNS_7 $T=2800 2490 0 0 $X=2700 $Y=2240
X15 6 7 4 8 6 pmos1v_CDNS_8 $T=4760 2040 0 0 $X=4340 $Y=1840
X16 8 7 4 nmos1v_CDNS_9 $T=4760 720 0 0 $X=4340 $Y=520
X17 6 5 1 8 6 pmos1v_CDNS_11 $T=930 2370 0 0 $X=510 $Y=2170
X18 8 5 1 nmos1v_CDNS_12 $T=930 850 0 0 $X=510 $Y=650
X19 8 5 9 8 nmos1v_CDNS_13 $T=2170 800 0 0 $X=1970 $Y=600
X20 4 3 10 8 nmos1v_CDNS_13 $T=3550 790 0 0 $X=3350 $Y=590
X21 4 2 9 8 nmos1v_CDNS_14 $T=1960 800 0 0 $X=1540 $Y=600
X22 8 1 10 8 nmos1v_CDNS_14 $T=3340 790 0 0 $X=2920 $Y=590
X23 6 1 11 8 6 pmos1v_CDNS_15 $T=2170 2100 0 0 $X=1970 $Y=1900
X24 4 3 12 8 6 pmos1v_CDNS_15 $T=3550 2030 0 0 $X=3350 $Y=1830
X25 4 2 11 8 6 pmos1v_CDNS_16 $T=1960 2100 0 0 $X=1540 $Y=1900
X26 6 5 12 8 6 pmos1v_CDNS_16 $T=3340 2030 0 0 $X=2920 $Y=1830
M0 9 2 4 8 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1960 $Y=800 $dt=0
M1 8 5 9 8 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=2170 $Y=800 $dt=0
M2 10 1 8 8 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3340 $Y=790 $dt=0
M3 4 3 10 8 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3550 $Y=790 $dt=0
M4 11 2 4 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8977 scb=0.0131425 scc=0.000918217 $X=1960 $Y=2100 $dt=1
M5 6 1 11 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=2170 $Y=2100 $dt=1
M6 12 5 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=3340 $Y=2030 $dt=1
M7 4 3 12 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=3550 $Y=2030 $dt=1
.ends MUX_2to1___2X_forph2p2
