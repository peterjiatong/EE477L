* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 4bit_CSA                                     *
* Netlisted  : Sun Nov  3 06:47:35 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR2_1X                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR2_1X A B vdd! gnd! OUT 6 7
*.DEVICECLIMB
** N=10 EP=7 FDC=10
M0 6 A gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=650 $Y=860 $dt=0
M1 7 B gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1580 $Y=860 $dt=0
M2 9 B gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=3020 $Y=860 $dt=0
M3 OUT 6 10 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=3950 $Y=860 $dt=0
M4 gnd! 7 10 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4880 $Y=860 $dt=0
M5 OUT A 9 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5810 $Y=860 $dt=0
M6 8 B vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3020 $Y=2500 $dt=1
M7 OUT 6 8 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=3950 $Y=2500 $dt=1
M8 OUT 7 8 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=4880 $Y=2500 $dt=1
M9 vdd! A 8 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.2959 scb=0.00764059 scc=8.89329e-05 $X=5810 $Y=2500 $dt=1
.ends XOR2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X in_a vdd! gnd! in_b out
** N=6 EP=5 FDC=4
M0 6 in_a gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=620 $Y=720 $dt=0
M1 out in_b 6 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=830 $Y=720 $dt=0
M2 out in_a vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=620 $Y=2080 $dt=1
M3 vdd! in_b out vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=21.6767 scb=0.0202328 scc=0.0021948 $X=1030 $Y=2080 $dt=1
.ends NAND2_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_2X                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_2X vdd! gnd! in_a in_b out
** N=6 EP=5 FDC=4
M0 6 in_a gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=7.2e-15 AS=1.68e-14 PD=3.6e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=2.45e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=620 $Y=710 $dt=0
M1 out in_b 6 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=7.2e-15 PD=5.2e-07 PS=3.6e-07 fw=1.2e-07 sa=2.45e-07 sb=1.4e-07 sca=7.31073 scb=0.00435535 scc=4.26584e-05 $X=830 $Y=710 $dt=0
M2 out in_a vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=15.9511 scb=0.0138709 scc=0.00113792 $X=620 $Y=2070 $dt=1
M3 vdd! in_b out vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=15.9511 scb=0.0138709 scc=0.00113792 $X=1030 $Y=2070 $dt=1
.ends NAND2_2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 1_bit_Full_Adder_ver1                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 1_bit_Full_Adder_ver1 A B Cin gnd! vdd! Cout S 11 12
*.DEVICECLIMB
** N=23 EP=9 FDC=34
X28 B vdd! gnd! A 10 NAND2_1X $T=8400 -10 0 0 $X=8400 $Y=0
X29 10 vdd! gnd! 9 Cout NAND2_1X $T=10400 -10 0 0 $X=10400 $Y=0
X30 vdd! gnd! 8 Cin 9 NAND2_2X $T=6400 0 0 0 $X=6400 $Y=0
X31 A B vdd! gnd! 8 11 12 XOR2_1X $T=0 0 0 0 $X=0 $Y=0
X32 Cin 8 vdd! gnd! S 13 14 XOR2_1X $T=12400 0 0 0 $X=12400 $Y=0
M0 13 Cin vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=13050 $Y=2490 $dt=1
M1 14 8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=13980 $Y=2490 $dt=1
.ends 1_bit_Full_Adder_ver1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X out vdd! gnd! in
** N=4 EP=4 FDC=2
M0 out in gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6908 scb=0.0179614 scc=0.00130074 $X=1090 $Y=1110 $dt=0
M1 out in vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=18.2452 scb=0.0177397 scc=0.00150411 $X=1090 $Y=2120 $dt=1
.ends INV_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND4_1x                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND4_1x B A vdd! gnd! C D OUT
** N=15 EP=7 FDC=18
X0 A vdd! gnd! B 8 NAND2_1X $T=0 -10 0 0 $X=0 $Y=0
X1 C vdd! gnd! D 9 NAND2_1X $T=4000 -10 0 0 $X=4000 $Y=0
X2 10 vdd! gnd! 11 12 NAND2_1X $T=8000 -10 0 0 $X=8000 $Y=0
X5 11 vdd! gnd! 8 INV_1X $T=1990 0 0 0 $X=2000 $Y=0
X6 10 vdd! gnd! 9 INV_1X $T=5990 0 0 0 $X=6000 $Y=0
X7 OUT vdd! gnd! 12 INV_1X $T=9990 0 0 0 $X=10000 $Y=0
.ends AND4_1x

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_1X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_1X vdd! S gnd! A B Out
** N=12 EP=6 FDC=12
M0 7 S gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=750 $Y=890 $dt=0
M1 9 7 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=2140 $Y=890 $dt=0
M2 11 S gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=3070 $Y=890 $dt=0
M3 8 A 9 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=4000 $Y=890 $dt=0
M4 8 B 11 gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=4930 $Y=890 $dt=0
M5 Out 8 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=6310 $Y=890 $dt=0
M6 7 S vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=750 $Y=2330 $dt=1
M7 10 7 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=2140 $Y=2330 $dt=1
M8 12 S vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=3070 $Y=2330 $dt=1
M9 8 A 12 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=4000 $Y=2330 $dt=1
M10 8 B 10 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=4930 $Y=2330 $dt=1
M11 Out 8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=19.0824 scb=0.0208702 scc=0.000619562 $X=6310 $Y=2330 $dt=1
.ends MUX_1X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 4bit_CSA                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 4bit_CSA A0 A1 A2 A3 B0 B1 B2 B3 C0 Cout
+ S0 S1 S2 S3 gnd! vdd!
** N=123 EP=16 FDC=222
X48 A0 B0 vdd! gnd! 5 26 27 XOR2_1X $T=18800 0 0 0 $X=18800 $Y=0
X49 A1 B1 vdd! gnd! 6 28 29 XOR2_1X $T=44000 0 0 0 $X=44000 $Y=0
X50 A2 B2 vdd! gnd! 7 30 31 XOR2_1X $T=69200 0 0 0 $X=69200 $Y=0
X51 A3 B3 vdd! gnd! 16 32 33 XOR2_1X $T=94400 0 0 0 $X=94400 $Y=0
X52 A0 B0 C0 gnd! vdd! 17 S0 34 35 1_bit_Full_Adder_ver1 $T=0 0 0 0 $X=0 $Y=0
X53 A1 B1 17 gnd! vdd! 19 S1 41 42 1_bit_Full_Adder_ver1 $T=25200 0 0 0 $X=25200 $Y=0
X54 A2 B2 19 gnd! vdd! 21 S2 48 49 1_bit_Full_Adder_ver1 $T=50400 0 0 0 $X=50400 $Y=0
X55 A3 B3 21 gnd! vdd! 12 S3 55 56 1_bit_Full_Adder_ver1 $T=75600 0 0 0 $X=75600 $Y=0
X56 7 16 vdd! gnd! 6 5 24 AND4_1x $T=100800 0 0 0 $X=100800 $Y=0
X57 vdd! 24 gnd! 12 C0 Cout MUX_1X $T=112790 0 0 0 $X=112800 $Y=0
M0 34 A0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=17.6861 scb=0.0184591 scc=0.000433664 $X=650 $Y=2490 $dt=1
M1 35 B0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.886 scb=0.00790338 scc=9.25552e-05 $X=1580 $Y=2490 $dt=1
M2 26 A0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=19450 $Y=2490 $dt=1
M3 27 B0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=20380 $Y=2490 $dt=1
M4 41 A1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=25850 $Y=2490 $dt=1
M5 42 B1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=26780 $Y=2490 $dt=1
M6 28 A1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=44650 $Y=2490 $dt=1
M7 29 B1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=45580 $Y=2490 $dt=1
M8 48 A2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=51050 $Y=2490 $dt=1
M9 49 B2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=51980 $Y=2490 $dt=1
M10 30 A2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=69850 $Y=2490 $dt=1
M11 31 B2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=70780 $Y=2490 $dt=1
M12 55 A3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=76250 $Y=2490 $dt=1
M13 56 B3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=77180 $Y=2490 $dt=1
M14 32 A3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=95050 $Y=2490 $dt=1
M15 33 B3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.327 scb=0.00769864 scc=9.24832e-05 $X=95980 $Y=2490 $dt=1
.ends 4bit_CSA
