* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : 10badder                                     *
* Netlisted  : Sun Nov 17 17:58:28 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X S gnd! vdd! A B out
** N=12 EP=6 FDC=12
M0 7 S gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=750 $Y=-4370 $dt=0
M1 9 A 8 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1780 $Y=-4420 $dt=0
M2 gnd! 7 9 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1990 $Y=-4420 $dt=0
M3 10 S gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3160 $Y=-4430 $dt=0
M4 8 B 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3370 $Y=-4430 $dt=0
M5 out 8 gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=4580 $Y=-4500 $dt=0
M6 7 S vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=750 $Y=-2850 $dt=1
M7 11 A 8 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1780 $Y=-3120 $dt=1
M8 vdd! S 11 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1990 $Y=-3120 $dt=1
M9 12 7 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3160 $Y=-3190 $dt=1
M10 8 B 12 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3370 $Y=-3190 $dt=1
M11 out 8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.2373 scb=0.0194294 scc=0.00149528 $X=4580 $Y=-3180 $dt=1
.ends MUX_2to1___2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_1X_small                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_1X_small vdd! gnd! 3 4 5
*.DEVICECLIMB
** N=6 EP=5 FDC=2
M0 6 3 gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1000 $Y=830 $dt=0
M1 4 5 6 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1210 $Y=830 $dt=0
.ends NAND_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR1 vdd! gnd! 3 4 5 6 7 9
*.DEVICECLIMB
** N=10 EP=8 FDC=6
M0 6 3 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=830 $Y=840 $dt=0
M1 7 4 gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1790 $Y=840 $dt=0
M2 8 4 gnd! gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=3120 $Y=780 $dt=0
M3 5 6 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4126 scb=0.0095497 scc=0.000351079 $X=4090 $Y=760 $dt=0
M4 gnd! 7 10 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=5050 $Y=770 $dt=0
M5 5 3 8 gnd! g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=6010 $Y=770 $dt=0
.ends XOR1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_2X_small1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_2X_small1 vdd! gnd! out 4 5
*.DEVICECLIMB
** N=6 EP=5 FDC=2
M0 6 4 gnd! gnd! g45n1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=7.66878 scb=0.00580736 scc=7.77234e-05 $X=940 $Y=890 $dt=0
M1 out 5 6 gnd! g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=11.676 scb=0.0124835 scc=0.000479408 $X=940 $Y=1100 $dt=0
.ends NAND_2X_small1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder1_small                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder1_small inA inB vdd! gnd! Cin_ S Cout 8 9 10
+ 11 12 13 14 22 23
*.DEVICECLIMB
** N=23 EP=16 FDC=18
X26 vdd! gnd! inA 10 inB NAND_1X_small $T=16970 30 0 0 $X=16540 $Y=10
X27 vdd! gnd! 9 Cout 10 NAND_1X_small $T=19810 30 0 0 $X=19380 $Y=10
X28 vdd! gnd! 9 Cin_ 8 NAND_2X_small1 $T=13690 -10 0 0 $X=13700 $Y=10
X29 vdd! gnd! inA inB 8 11 12 22 XOR1 $T=-40 30 0 0 $X=20 $Y=10
X30 vdd! gnd! Cin_ 8 S 13 14 23 XOR1 $T=6800 30 0 0 $X=6860 $Y=10
.ends full_adder1_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FA_4bit                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FA_4bit vdd! B0 A0 B1 A1 B2 A2 B3 A3 gnd!
+ Cin_rrr S0 S1 S2 S3 Cout3
** N=83 EP=16 FDC=144
X20 A0 B0 vdd! gnd! Cin_rrr S0 17 43 46 47
+ 41 42 44 45 82 83 full_adder1_small $T=-90 -130 0 0 $X=-70 $Y=-120
X21 A1 B1 vdd! gnd! 17 S1 19 36 39 40
+ 34 35 37 38 80 81 full_adder1_small $T=-90 7250 1 0 $X=-70 $Y=3440
X22 A2 B2 vdd! gnd! 19 S2 18 29 32 33
+ 27 28 30 31 78 79 full_adder1_small $T=-90 7190 0 0 $X=-70 $Y=7200
X23 A3 B3 vdd! gnd! 18 S3 Cout3 22 25 26
+ 20 21 23 24 76 77 full_adder1_small $T=-90 14570 1 0 $X=-70 $Y=10760
M0 41 A0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=2220 $dt=1
M1 34 A1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=4420 $dt=1
M2 27 A2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=9540 $dt=1
M3 20 A3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=11740 $dt=1
M4 42 B0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=2220 $dt=1
M5 35 B1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=4420 $dt=1
M6 28 B2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=9540 $dt=1
M7 21 B3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=11740 $dt=1
M8 82 B0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=1980 $dt=1
M9 80 B1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=4180 $dt=1
M10 78 B2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=9300 $dt=1
M11 76 B3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=11500 $dt=1
M12 43 41 82 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=2040 $dt=1
M13 36 34 80 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=4120 $dt=1
M14 29 27 78 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=9360 $dt=1
M15 22 20 76 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=11440 $dt=1
M16 43 42 82 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=2040 $dt=1
M17 36 35 80 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=4120 $dt=1
M18 29 28 78 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=9360 $dt=1
M19 22 21 76 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=11440 $dt=1
M20 82 A0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=2040 $dt=1
M21 80 A1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=4120 $dt=1
M22 78 A2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=9360 $dt=1
M23 76 A3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=11440 $dt=1
M24 44 Cin_rrr vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=2220 $dt=1
M25 37 17 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=4420 $dt=1
M26 30 19 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=9540 $dt=1
M27 23 18 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=11740 $dt=1
M28 45 43 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=2220 $dt=1
M29 38 36 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=4420 $dt=1
M30 31 29 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=9540 $dt=1
M31 24 22 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=11740 $dt=1
M32 83 43 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=1980 $dt=1
M33 81 36 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=4180 $dt=1
M34 79 29 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=9300 $dt=1
M35 77 22 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=11500 $dt=1
M36 S0 44 83 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=2040 $dt=1
M37 S1 37 81 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=4120 $dt=1
M38 S2 30 79 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=9360 $dt=1
M39 S3 23 77 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=11440 $dt=1
M40 S0 45 83 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=2040 $dt=1
M41 S1 38 81 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=4120 $dt=1
M42 S2 31 79 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=9360 $dt=1
M43 S3 24 77 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=11440 $dt=1
M44 83 Cin_rrr vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=2040 $dt=1
M45 81 17 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=4120 $dt=1
M46 79 19 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=9360 $dt=1
M47 77 18 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=11440 $dt=1
M48 46 Cin_rrr vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=2010 $dt=1
M49 39 17 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=4150 $dt=1
M50 32 19 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=9330 $dt=1
M51 25 18 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=11470 $dt=1
M52 vdd! 43 46 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=2010 $dt=1
M53 vdd! 36 39 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=4150 $dt=1
M54 vdd! 29 32 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=9330 $dt=1
M55 vdd! 22 25 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=11470 $dt=1
M56 47 A0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=2230 $dt=1
M57 40 A1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=4410 $dt=1
M58 33 A2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=9550 $dt=1
M59 26 A3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=11730 $dt=1
M60 vdd! B0 47 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=2230 $dt=1
M61 vdd! B1 40 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=4410 $dt=1
M62 vdd! B2 33 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=9550 $dt=1
M63 vdd! B3 26 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=11730 $dt=1
M64 17 46 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=2230 $dt=1
M65 19 39 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=4410 $dt=1
M66 18 32 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=9550 $dt=1
M67 Cout3 25 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=11730 $dt=1
M68 vdd! 47 17 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=2230 $dt=1
M69 vdd! 40 19 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=4410 $dt=1
M70 vdd! 33 18 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=9550 $dt=1
M71 vdd! 26 Cout3 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=11730 $dt=1
.ends FA_4bit

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small in vdd! gnd! out
** N=4 EP=4 FDC=2
M0 out in gnd! gnd! g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7353 scb=0.0117274 scc=0.000445561 $X=1070 $Y=980 $dt=0
M1 out in vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8675 scb=0.0146094 scc=0.000688105 $X=1070 $Y=2220 $dt=1
.ends INV_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 10badder                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 10badder Cin Cout S0 S1 S2 S3 S4 S5 S6 S7
+ S8 S9 gnd! in_A_0 in_A_1 in_A_2 in_A_3 in_A_4 in_A_5 in_A_6
+ in_A_7 in_A_8 in_A_9 in_B_0 in_B_1 in_B_2 in_B_3 in_B_4 in_B_5 in_B_6
+ in_B_7 in_B_8 in_B_9 vdd!
** N=267 EP=34 FDC=516
X147 26 gnd! vdd! 2 Cin 1 MUX_2to1___2X $T=56190 30160 0 180 $X=50640 $Y=31580
X148 27 gnd! vdd! 3 1 4 MUX_2to1___2X $T=56190 44800 0 180 $X=50640 $Y=46220
X149 vdd! gnd! 11 34 13 NAND_1X_small $T=53960 20720 0 0 $X=53530 $Y=20700
X150 vdd! gnd! 9 36 28 NAND_1X_small $T=55940 28040 0 180 $X=53530 $Y=24260
X151 vdd! gnd! 7 32 15 NAND_1X_small $T=53960 28040 0 0 $X=53530 $Y=28020
X152 vdd! gnd! 12 35 14 NAND_1X_small $T=53960 35360 0 0 $X=53530 $Y=35340
X153 vdd! gnd! 10 37 29 NAND_1X_small $T=55940 42680 0 180 $X=53530 $Y=38900
X154 vdd! gnd! 8 33 16 NAND_1X_small $T=53960 42680 0 0 $X=53530 $Y=42660
X155 vdd! gnd! in_B_0 in_A_0 13 64 65 256 XOR1 $T=56070 20720 0 0 $X=56130 $Y=20700
X156 vdd! gnd! in_A_1 in_B_1 11 66 67 257 XOR1 $T=56070 28040 1 0 $X=56130 $Y=24260
X157 vdd! gnd! in_A_2 in_B_2 15 68 69 258 XOR1 $T=56070 28040 0 0 $X=56130 $Y=28020
X158 vdd! gnd! in_A_3 in_B_3 7 70 71 259 XOR1 $T=56070 35360 1 0 $X=56130 $Y=31580
X159 vdd! gnd! in_B_4 in_A_4 14 72 73 260 XOR1 $T=56070 35360 0 0 $X=56130 $Y=35340
X160 vdd! gnd! in_A_5 in_B_5 12 74 75 261 XOR1 $T=56070 42680 1 0 $X=56130 $Y=38900
X161 vdd! gnd! in_A_6 in_B_6 16 76 77 262 XOR1 $T=56070 42680 0 0 $X=56130 $Y=42660
X162 vdd! gnd! in_A_7 in_B_7 8 78 79 263 XOR1 $T=56070 50000 1 0 $X=56130 $Y=46220
X163 in_B_8 in_A_8 vdd! gnd! 4 S8 5 82 85 86
+ 80 81 83 84 264 265 full_adder1_small $T=50650 49970 0 0 $X=50670 $Y=49980
X164 in_A_9 in_B_9 vdd! gnd! 5 S9 Cout 89 92 93
+ 87 88 90 91 266 267 full_adder1_small $T=72610 49970 0 0 $X=72630 $Y=49980
X165 vdd! in_B_0 in_A_0 in_B_1 in_A_1 in_B_2 in_A_2 in_B_3 in_A_3 gnd!
+ Cin S0 S1 S2 S3 2 FA_4bit $T=64900 20820 0 0 $X=64250 $Y=20700
X166 vdd! in_B_4 in_A_4 in_B_5 in_A_5 in_B_6 in_A_6 in_B_7 in_A_7 gnd!
+ 1 S4 S5 S6 S7 3 FA_4bit $T=64900 35460 0 0 $X=64250 $Y=35340
X167 34 vdd! gnd! 28 INV_1X_small $T=51530 20700 0 0 $X=51530 $Y=20700
X168 36 vdd! gnd! 26 INV_1X_small $T=51530 28060 1 0 $X=51530 $Y=24260
X169 32 vdd! gnd! 9 INV_1X_small $T=51530 28020 0 0 $X=51530 $Y=28020
X170 35 vdd! gnd! 29 INV_1X_small $T=51530 35340 0 0 $X=51530 $Y=35340
X171 37 vdd! gnd! 27 INV_1X_small $T=51530 42700 1 0 $X=51530 $Y=38900
X172 33 vdd! gnd! 10 INV_1X_small $T=51530 42660 0 0 $X=51530 $Y=42660
M0 80 in_B_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6612 scb=0.0167915 scc=0.000377457 $X=51440 $Y=52320 $dt=1
M1 81 in_A_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.8911 scb=0.00996238 scc=0.000256798 $X=52400 $Y=52320 $dt=1
M2 264 in_A_8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=53730 $Y=52080 $dt=1
M3 36 28 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=25230 $dt=1
M4 37 29 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=39870 $dt=1
M5 82 80 264 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=54700 $Y=52140 $dt=1
M6 34 11 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=23050 $dt=1
M7 32 7 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=30370 $dt=1
M8 35 12 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=37690 $dt=1
M9 33 8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=45010 $dt=1
M10 vdd! 9 36 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=25230 $dt=1
M11 vdd! 10 37 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=39870 $dt=1
M12 vdd! 13 34 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=23050 $dt=1
M13 vdd! 15 32 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=30370 $dt=1
M14 vdd! 14 35 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=37690 $dt=1
M15 vdd! 16 33 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=45010 $dt=1
M16 82 81 264 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=55660 $Y=52140 $dt=1
M17 264 in_B_8 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=56620 $Y=52140 $dt=1
M18 64 in_B_0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=23040 $dt=1
M19 66 in_A_1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=25240 $dt=1
M20 68 in_A_2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=30360 $dt=1
M21 70 in_A_3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=32560 $dt=1
M22 72 in_B_4 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=37680 $dt=1
M23 74 in_A_5 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=39880 $dt=1
M24 76 in_A_6 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=45000 $dt=1
M25 78 in_A_7 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=47200 $dt=1
M26 65 in_A_0 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=23040 $dt=1
M27 67 in_B_1 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=25240 $dt=1
M28 69 in_B_2 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=30360 $dt=1
M29 71 in_B_3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=32560 $dt=1
M30 73 in_A_4 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=37680 $dt=1
M31 75 in_B_5 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=39880 $dt=1
M32 77 in_B_6 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=45000 $dt=1
M33 79 in_B_7 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=47200 $dt=1
M34 83 4 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=58280 $Y=52320 $dt=1
M35 256 in_A_0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=22800 $dt=1
M36 257 in_B_1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=25000 $dt=1
M37 258 in_B_2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=30120 $dt=1
M38 259 in_B_3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=32320 $dt=1
M39 260 in_A_4 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=37440 $dt=1
M40 261 in_B_5 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=39640 $dt=1
M41 262 in_B_6 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=44760 $dt=1
M42 263 in_B_7 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=46960 $dt=1
M43 84 82 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=59240 $Y=52320 $dt=1
M44 13 64 256 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=22860 $dt=1
M45 11 66 257 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=24940 $dt=1
M46 15 68 258 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=30180 $dt=1
M47 7 70 259 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=32260 $dt=1
M48 14 72 260 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=37500 $dt=1
M49 12 74 261 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=39580 $dt=1
M50 16 76 262 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=44820 $dt=1
M51 8 78 263 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=46900 $dt=1
M52 265 82 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60570 $Y=52080 $dt=1
M53 13 65 256 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=22860 $dt=1
M54 11 67 257 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=24940 $dt=1
M55 15 69 258 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=30180 $dt=1
M56 7 71 259 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=32260 $dt=1
M57 14 73 260 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=37500 $dt=1
M58 12 75 261 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=39580 $dt=1
M59 16 77 262 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=44820 $dt=1
M60 8 79 263 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=46900 $dt=1
M61 S8 83 265 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=61540 $Y=52140 $dt=1
M62 256 in_B_0 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=22860 $dt=1
M63 257 in_A_1 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=24940 $dt=1
M64 258 in_A_2 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=30180 $dt=1
M65 259 in_A_3 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=32260 $dt=1
M66 260 in_B_4 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=37500 $dt=1
M67 261 in_A_5 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=39580 $dt=1
M68 262 in_A_6 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=44820 $dt=1
M69 263 in_A_7 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=46900 $dt=1
M70 S8 84 265 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=62500 $Y=52140 $dt=1
M71 265 4 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=63460 $Y=52140 $dt=1
M72 85 4 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65530 $Y=52110 $dt=1
M73 vdd! 82 85 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65940 $Y=52110 $dt=1
M74 86 in_B_8 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68510 $Y=52330 $dt=1
M75 vdd! in_A_8 86 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68920 $Y=52330 $dt=1
M76 5 85 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71350 $Y=52330 $dt=1
M77 vdd! 86 5 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71760 $Y=52330 $dt=1
M78 87 in_A_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=73400 $Y=52320 $dt=1
M79 88 in_B_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=74360 $Y=52320 $dt=1
M80 266 in_B_9 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=75690 $Y=52080 $dt=1
M81 89 87 266 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=76660 $Y=52140 $dt=1
M82 89 88 266 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=77620 $Y=52140 $dt=1
M83 266 in_A_9 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=78580 $Y=52140 $dt=1
M84 90 5 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=80240 $Y=52320 $dt=1
M85 91 89 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=81200 $Y=52320 $dt=1
M86 267 89 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=82530 $Y=52080 $dt=1
M87 S9 90 267 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=83500 $Y=52140 $dt=1
M88 S9 91 267 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=84460 $Y=52140 $dt=1
M89 267 5 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=85420 $Y=52140 $dt=1
M90 92 5 vdd! vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87490 $Y=52110 $dt=1
M91 vdd! 89 92 vdd! g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87900 $Y=52110 $dt=1
M92 93 in_A_9 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90470 $Y=52330 $dt=1
M93 vdd! in_B_9 93 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90880 $Y=52330 $dt=1
M94 Cout 92 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=93310 $Y=52330 $dt=1
M95 vdd! 93 Cout vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=93720 $Y=52330 $dt=1
.ends 10badder
