* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : OR2_1X                                       *
* Netlisted  : Wed Nov  6 21:04:10 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_4 D_drain_1 S_source_0 3
** N=3 EP=3 FDC=1
M0 D_drain_1 3 S_source_0 S_source_0 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: OR2_1X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt OR2_1X gnd! in_A in_B out vdd!
** N=7 EP=5 FDC=6
X6 3 gnd! in_A nmos1v_CDNS_4 $T=740 890 0 0 $X=320 $Y=690
X7 3 gnd! in_B nmos1v_CDNS_4 $T=1670 890 0 0 $X=1250 $Y=690
X8 out gnd! 3 nmos1v_CDNS_4 $T=2600 890 0 0 $X=2180 $Y=690
M0 4 in_A vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.75 scb=0.0169824 scc=0.000359091 $X=740 $Y=2370 $dt=1
M1 3 in_B 4 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.9866 scb=0.00948303 scc=0.000202299 $X=1670 $Y=2370 $dt=1
M2 out 3 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.5867 scb=0.0166976 scc=0.000345988 $X=2600 $Y=2370 $dt=1
.ends OR2_1X
