* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph2p2_processing_element                     *
* Netlisted  : Sun Nov 24 19:46:07 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_8                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_8 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_9                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_9 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_10                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_10 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_11                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_11 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_12                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_12 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_13                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_13 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_14                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_14 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_15                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_15 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_16                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_16 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_17                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_17 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_18                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_18 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_new                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_new 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 3 M1_PO_CDNS_16 $T=1020 1750 0 90 $X=900 $Y=1650
X1 1 2 cellTmpl_CDNS_18 $T=50 150 0 0 $X=-70 $Y=10
M0 4 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.3086 scb=0.00950139 scc=0.000267597 $X=1140 $Y=930 $dt=0
.ends INV_1X_new

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_19                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_19 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_20                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_20 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_20

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_21                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_21 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_21

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X_small                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_16 $T=690 1680 0 90 $X=570 $Y=1580
X1 4 M1_PO_CDNS_16 $T=1930 1650 0 90 $X=1810 $Y=1550
X2 3 1 6 3 nmos1v_CDNS_19 $T=810 1000 0 0 $X=390 $Y=800
X3 6 4 5 3 nmos1v_CDNS_19 $T=2050 1000 0 0 $X=1630 $Y=800
X4 2 1 5 3 2 pmos1v_CDNS_20 $T=810 2440 0 0 $X=390 $Y=2240
X5 2 4 5 3 2 pmos1v_CDNS_20 $T=2050 2450 0 0 $X=1630 $Y=2250
X6 2 3 cellTmpl_CDNS_21 $T=240 210 0 0 $X=120 $Y=70
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=810 $Y=1000 $dt=0
M1 5 4 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=2050 $Y=1000 $dt=0
.ends NAND2_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6
*.DEVICECLIMB
** N=7 EP=6 FDC=3
X0 2 3 6 5 INV_1X_new $T=2480 -10 0 0 $X=2410 $Y=0
X1 1 2 3 4 6 7 NAND2_1X_small $T=-110 -70 0 0 $X=10 $Y=0
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_22                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_22 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_23                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_23 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_23

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_24                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_24 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_24

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_25                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_25 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_25

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_26                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_26 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_26

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_27                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_27 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_27

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_28                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_28 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_28

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_29                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_29 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_29

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR_small                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR_small 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=9
X0 1 M2_M1_CDNS_8 $T=350 1340 0 90 $X=220 $Y=1260
X1 6 M2_M1_CDNS_8 $T=5510 3180 0 90 $X=5380 $Y=3100
X2 6 M2_M1_CDNS_8 $T=6740 3180 0 90 $X=6610 $Y=3100
X3 1 M1_PO_CDNS_16 $T=580 1660 0 90 $X=460 $Y=1560
X4 4 M1_PO_CDNS_16 $T=1990 1480 0 90 $X=1870 $Y=1380
X5 4 M1_PO_CDNS_22 $T=5990 1680 0 90 $X=5790 $Y=1580
X6 1 M1_PO_CDNS_22 $T=7100 1350 0 90 $X=6900 $Y=1250
X7 7 M1_PO_CDNS_23 $T=3070 1660 0 90 $X=2870 $Y=1560
X8 8 M1_PO_CDNS_23 $T=4410 1540 0 90 $X=4210 $Y=1440
X9 8 M3_M2_CDNS_24 $T=1210 1540 0 90 $X=1010 $Y=1440
X10 8 M3_M2_CDNS_24 $T=4410 1540 0 90 $X=4210 $Y=1440
X11 8 M2_M1_CDNS_25 $T=1210 1540 0 90 $X=1010 $Y=1440
X12 4 M2_M1_CDNS_25 $T=1820 1880 0 90 $X=1620 $Y=1780
X13 8 M2_M1_CDNS_25 $T=4410 1540 0 90 $X=4210 $Y=1440
X14 4 M2_M1_CDNS_26 $T=5990 1680 0 90 $X=5790 $Y=1580
X15 1 M2_M1_CDNS_26 $T=7100 1350 0 90 $X=6900 $Y=1250
X16 2 3 cellTmpl_CDNS_27 $T=120 140 0 0 $X=0 $Y=0
X17 2 1 8 3 2 pmos1v_CDNS_28 $T=700 2180 0 0 $X=280 $Y=1980
X18 2 4 7 3 2 pmos1v_CDNS_28 $T=2110 2170 0 0 $X=1690 $Y=1970
X19 2 7 6 3 2 pmos1v_CDNS_28 $T=3270 2160 0 0 $X=2850 $Y=1960
X20 2 8 6 3 2 pmos1v_CDNS_28 $T=4610 2160 0 0 $X=4190 $Y=1960
X21 6 4 5 3 2 pmos1v_CDNS_28 $T=6140 2120 0 0 $X=5720 $Y=1920
X22 6 1 5 3 2 pmos1v_CDNS_28 $T=7250 2160 0 0 $X=6830 $Y=1960
X23 3 1 8 3 nmos1v_CDNS_29 $T=700 590 0 0 $X=280 $Y=390
X24 3 4 7 3 nmos1v_CDNS_29 $T=2110 580 0 0 $X=1690 $Y=380
X25 3 7 9 3 nmos1v_CDNS_29 $T=3270 580 0 0 $X=2850 $Y=380
X26 9 8 5 3 nmos1v_CDNS_29 $T=4610 580 0 0 $X=4190 $Y=380
X27 3 4 10 3 nmos1v_CDNS_29 $T=6140 600 0 0 $X=5720 $Y=400
X28 10 1 5 3 nmos1v_CDNS_29 $T=7250 650 0 0 $X=6830 $Y=450
M0 8 1 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.45462 scb=0.00478425 scc=6.8709e-05 $X=700 $Y=590 $dt=0
M1 7 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=2110 $Y=580 $dt=0
M2 9 7 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=3270 $Y=580 $dt=0
M3 5 8 9 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=4610 $Y=580 $dt=0
M4 10 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 $X=6140 $Y=600 $dt=0
M5 5 1 10 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=7250 $Y=650 $dt=0
M6 7 4 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.1869 scb=0.0086398 scc=0.00051649 $X=2110 $Y=2170 $dt=1
M7 6 7 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3270 $Y=2160 $dt=1
M8 6 8 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4610 $Y=2160 $dt=1
.ends XOR_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 8 9 13
*.DEVICECLIMB
** N=13 EP=9 FDC=12
X0 4 M2_M1_CDNS_3 $T=6750 2480 0 0 $X=6670 $Y=2230
X1 4 M2_M1_CDNS_3 $T=9120 2880 0 0 $X=9040 $Y=2630
X2 4 M1_PO_CDNS_6 $T=6750 2480 0 0 $X=6650 $Y=2230
X3 4 M1_PO_CDNS_6 $T=9120 2880 0 0 $X=9020 $Y=2630
X4 4 M3_M2_CDNS_9 $T=6750 2480 0 0 $X=6670 $Y=2230
X5 4 M3_M2_CDNS_9 $T=9120 2880 0 0 $X=9040 $Y=2630
X6 1 3 2 4 6 9 AND $T=7790 0 0 0 $X=7800 $Y=0
X7 1 3 2 4 5 13 7 8 10 11 XOR_small $T=0 0 0 0 $X=0 $Y=0
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_33                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_33 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_33

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_1X_small                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=-310 120 0 0 $X=-430 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1000 $Y=830 $dt=0
M1 4 5 6 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1210 $Y=830 $dt=0
.ends NAND_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_2X_small1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_2X_small1 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=130 160 0 0 $X=10 $Y=20
M0 6 4 2 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=7.66878 scb=0.00580736 scc=7.77234e-05 $X=940 $Y=890 $dt=0
M1 3 5 6 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=11.676 scb=0.0124835 scc=0.000479408 $X=940 $Y=1100 $dt=0
.ends NAND_2X_small1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_39                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_39 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_39

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR1 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=6
X0 6 M2_M1_CDNS_8 $T=1210 1480 0 90 $X=1080 $Y=1400
X1 7 M2_M1_CDNS_8 $T=2250 1860 0 90 $X=2120 $Y=1780
X2 6 M2_M1_CDNS_8 $T=2950 1480 0 90 $X=2820 $Y=1400
X3 8 M2_M1_CDNS_8 $T=3370 650 0 0 $X=3290 $Y=520
X4 9 M2_M1_CDNS_8 $T=3370 3080 0 0 $X=3290 $Y=2950
X5 9 M2_M1_CDNS_8 $T=3930 3080 0 0 $X=3850 $Y=2950
X6 7 M2_M1_CDNS_8 $T=4680 1860 0 90 $X=4550 $Y=1780
X7 9 M2_M1_CDNS_8 $T=4890 3070 0 0 $X=4810 $Y=2940
X8 8 M2_M1_CDNS_8 $T=5840 640 0 0 $X=5760 $Y=510
X9 9 M2_M1_CDNS_8 $T=6260 3080 0 0 $X=6180 $Y=2950
X10 6 M1_PO_CDNS_16 $T=4020 1500 0 90 $X=3900 $Y=1400
X11 7 M1_PO_CDNS_16 $T=5020 1730 0 90 $X=4900 $Y=1630
X12 2 3 6 2 nmos1v_CDNS_19 $T=830 840 0 0 $X=410 $Y=640
X13 2 4 7 2 nmos1v_CDNS_19 $T=1790 840 0 0 $X=1370 $Y=640
X14 1 3 6 2 1 pmos1v_CDNS_20 $T=830 2320 0 0 $X=410 $Y=2120
X15 1 4 7 2 1 pmos1v_CDNS_20 $T=1790 2320 0 0 $X=1370 $Y=2120
X16 1 4 9 2 1 pmos1v_CDNS_28 $T=3120 2080 0 0 $X=2700 $Y=1880
X17 9 6 5 2 1 pmos1v_CDNS_28 $T=4090 2140 0 0 $X=3670 $Y=1940
X18 9 7 5 2 1 pmos1v_CDNS_28 $T=5050 2140 0 0 $X=4630 $Y=1940
X19 1 3 9 2 1 pmos1v_CDNS_28 $T=6010 2140 0 0 $X=5590 $Y=1940
X20 2 4 8 2 nmos1v_CDNS_29 $T=3120 780 0 0 $X=2700 $Y=580
X21 10 6 5 2 nmos1v_CDNS_29 $T=4090 760 0 0 $X=3670 $Y=560
X22 10 7 2 2 nmos1v_CDNS_29 $T=5050 770 0 0 $X=4630 $Y=570
X23 8 3 5 2 nmos1v_CDNS_29 $T=6010 770 0 0 $X=5590 $Y=570
X24 1 2 cellTmpl_CDNS_39 $T=180 120 0 0 $X=60 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=830 $Y=840 $dt=0
M1 7 4 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1790 $Y=840 $dt=0
M2 8 4 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=3120 $Y=780 $dt=0
M3 5 6 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4126 scb=0.0095497 scc=0.000351079 $X=4090 $Y=760 $dt=0
M4 2 7 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=5050 $Y=770 $dt=0
M5 5 3 8 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=6010 $Y=770 $dt=0
.ends XOR1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder1_small                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder1_small 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 22 23
*.DEVICECLIMB
** N=23 EP=16 FDC=18
X0 1 M2_M1_CDNS_3 $T=590 2080 0 90 $X=340 $Y=2000
X1 3 M2_M1_CDNS_3 $T=2300 3150 0 90 $X=2050 $Y=3070
X2 1 M2_M1_CDNS_3 $T=17380 1890 0 0 $X=17300 $Y=1640
X3 3 M2_M1_CDNS_3 $T=19040 3010 0 0 $X=18960 $Y=2760
X4 1 M1_PO_CDNS_6 $T=590 2080 0 90 $X=340 $Y=1980
X5 3 M1_PO_CDNS_6 $T=2300 3150 0 90 $X=2050 $Y=3050
X6 1 M1_PO_CDNS_6 $T=17380 1890 0 0 $X=17280 $Y=1640
X7 3 M1_PO_CDNS_6 $T=19040 3010 0 0 $X=18940 $Y=2760
X8 8 M2_M1_CDNS_8 $T=6580 1900 0 0 $X=6500 $Y=1770
X9 9 M2_M1_CDNS_8 $T=15190 1730 0 90 $X=15060 $Y=1650
X10 1 M3_M2_CDNS_9 $T=590 2080 0 90 $X=340 $Y=2000
X11 3 M3_M2_CDNS_9 $T=2300 3150 0 90 $X=2050 $Y=3070
X12 1 M3_M2_CDNS_9 $T=17380 1890 0 0 $X=17300 $Y=1640
X13 3 M3_M2_CDNS_9 $T=19040 3010 0 0 $X=18960 $Y=2760
X14 8 M3_M2_CDNS_10 $T=6970 950 0 0 $X=6890 $Y=820
X15 8 M3_M2_CDNS_10 $T=14100 570 0 90 $X=13970 $Y=490
X16 8 M1_PO_CDNS_15 $T=8510 1970 0 0 $X=8410 $Y=1720
X17 8 M1_PO_CDNS_15 $T=16110 1570 0 0 $X=16010 $Y=1320
X18 9 M1_PO_CDNS_15 $T=20260 1840 0 0 $X=20160 $Y=1590
X19 1 M1_PO_CDNS_16 $T=690 1610 0 0 $X=590 $Y=1490
X20 3 M1_PO_CDNS_16 $T=1650 1990 0 0 $X=1550 $Y=1870
X21 5 M1_PO_CDNS_16 $T=7590 1960 0 0 $X=7490 $Y=1840
X22 10 M1_PO_CDNS_16 $T=19320 1680 0 0 $X=19220 $Y=1560
X23 8 M2_M1_CDNS_17 $T=8510 1970 0 0 $X=8430 $Y=1720
X24 8 M2_M1_CDNS_17 $T=16110 1570 0 0 $X=16030 $Y=1320
X25 9 M2_M1_CDNS_17 $T=20260 1840 0 0 $X=20180 $Y=1590
X26 2 4 1 10 3 20 NAND_1X_small $T=16970 30 0 0 $X=16540 $Y=10
X27 2 4 9 7 10 21 NAND_1X_small $T=19810 30 0 0 $X=19380 $Y=10
X28 2 4 9 5 8 19 NAND_2X_small1 $T=13690 -10 0 0 $X=13700 $Y=10
X29 2 4 1 3 8 11 12 15 22 16 XOR1 $T=-40 30 0 0 $X=20 $Y=10
X30 2 4 5 8 6 13 14 17 23 18 XOR1 $T=6800 30 0 0 $X=6860 $Y=10
.ends full_adder1_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: multiplier                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt multiplier 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
** N=238 EP=50 FDC=456
X0 1 M4_M3_CDNS_1 $T=1390 19500 0 0 $X=1310 $Y=19250
X1 19 M4_M3_CDNS_1 $T=3370 8280 0 0 $X=3290 $Y=8030
X2 7 M4_M3_CDNS_1 $T=4510 16920 0 0 $X=4430 $Y=16670
X3 20 M4_M3_CDNS_1 $T=5400 9800 0 0 $X=5320 $Y=9550
X4 7 M4_M3_CDNS_1 $T=7950 19550 0 0 $X=7870 $Y=19300
X5 21 M4_M3_CDNS_1 $T=8750 8160 0 0 $X=8670 $Y=7910
X6 22 M4_M3_CDNS_1 $T=10750 19470 0 0 $X=10670 $Y=19220
X7 23 M4_M3_CDNS_1 $T=11680 11800 0 0 $X=11600 $Y=11550
X8 24 M4_M3_CDNS_1 $T=12950 9830 0 0 $X=12870 $Y=9580
X9 11 M4_M3_CDNS_1 $T=13290 16990 0 0 $X=13210 $Y=16740
X10 25 M4_M3_CDNS_1 $T=14070 2580 0 90 $X=13820 $Y=2500
X11 26 M4_M3_CDNS_1 $T=15700 9710 0 0 $X=15620 $Y=9460
X12 23 M4_M3_CDNS_1 $T=22150 6400 0 0 $X=22070 $Y=6150
X13 26 M4_M3_CDNS_1 $T=24490 750 0 0 $X=24410 $Y=500
X14 11 M4_M3_CDNS_1 $T=25590 19380 0 0 $X=25510 $Y=19130
X15 27 M4_M3_CDNS_1 $T=25970 20660 0 0 $X=25890 $Y=20410
X16 28 M4_M3_CDNS_1 $T=26370 19410 0 0 $X=26290 $Y=19160
X17 29 M4_M3_CDNS_1 $T=26600 23000 0 0 $X=26520 $Y=22750
X18 30 M4_M3_CDNS_1 $T=28540 8430 0 0 $X=28460 $Y=8180
X19 30 M4_M3_CDNS_1 $T=28700 9810 0 0 $X=28620 $Y=9560
X20 31 M4_M3_CDNS_1 $T=29280 19170 0 0 $X=29200 $Y=18920
X21 32 M4_M3_CDNS_1 $T=35970 2380 0 0 $X=35890 $Y=2130
X22 33 M4_M3_CDNS_1 $T=38260 18710 0 0 $X=38180 $Y=18460
X23 31 M4_M3_CDNS_1 $T=39640 17490 0 0 $X=39560 $Y=17240
X24 32 M4_M3_CDNS_1 $T=42090 2930 0 90 $X=41840 $Y=2850
X25 34 M4_M3_CDNS_1 $T=43850 8260 0 0 $X=43770 $Y=8010
X26 35 M4_M3_CDNS_1 $T=43880 660 0 0 $X=43800 $Y=410
X27 33 M4_M3_CDNS_1 $T=46340 18970 0 0 $X=46260 $Y=18720
X28 1 M3_M2_CDNS_2 $T=1390 21140 0 0 $X=1310 $Y=20890
X29 7 M3_M2_CDNS_2 $T=4510 16920 0 0 $X=4430 $Y=16670
X30 21 M3_M2_CDNS_2 $T=8750 8160 0 0 $X=8670 $Y=7910
X31 22 M3_M2_CDNS_2 $T=10750 19470 0 0 $X=10670 $Y=19220
X32 23 M3_M2_CDNS_2 $T=11680 11800 0 0 $X=11600 $Y=11550
X33 27 M3_M2_CDNS_2 $T=13170 22790 0 0 $X=13090 $Y=22540
X34 11 M3_M2_CDNS_2 $T=13290 16990 0 0 $X=13210 $Y=16740
X35 11 M3_M2_CDNS_2 $T=14530 13310 0 0 $X=14450 $Y=13060
X36 11 M3_M2_CDNS_2 $T=14530 15600 0 0 $X=14450 $Y=15350
X37 23 M3_M2_CDNS_2 $T=22150 6400 0 0 $X=22070 $Y=6150
X38 26 M3_M2_CDNS_2 $T=24490 750 0 0 $X=24410 $Y=500
X39 28 M3_M2_CDNS_2 $T=26370 19410 0 0 $X=26290 $Y=19160
X40 29 M3_M2_CDNS_2 $T=26600 23000 0 0 $X=26520 $Y=22750
X41 36 M3_M2_CDNS_2 $T=28820 19250 0 0 $X=28740 $Y=19000
X42 31 M3_M2_CDNS_2 $T=29280 19170 0 0 $X=29200 $Y=18920
X43 22 M3_M2_CDNS_2 $T=33860 19960 0 90 $X=33610 $Y=19880
X44 36 M3_M2_CDNS_2 $T=34220 19150 0 0 $X=34140 $Y=18900
X45 32 M3_M2_CDNS_2 $T=35970 2380 0 0 $X=35890 $Y=2130
X46 31 M3_M2_CDNS_2 $T=39640 17490 0 0 $X=39560 $Y=17240
X47 34 M3_M2_CDNS_2 $T=43850 8260 0 0 $X=43770 $Y=8010
X48 35 M3_M2_CDNS_2 $T=43880 660 0 0 $X=43800 $Y=410
X49 33 M3_M2_CDNS_2 $T=46340 18970 0 0 $X=46260 $Y=18720
X50 1 M2_M1_CDNS_3 $T=1350 15570 0 0 $X=1270 $Y=15320
X51 1 M2_M1_CDNS_3 $T=1360 13320 0 0 $X=1280 $Y=13070
X52 1 M2_M1_CDNS_3 $T=1390 21140 0 0 $X=1310 $Y=20890
X53 7 M2_M1_CDNS_3 $T=4510 16920 0 0 $X=4430 $Y=16670
X54 7 M2_M1_CDNS_3 $T=5740 15570 0 0 $X=5660 $Y=15320
X55 7 M2_M1_CDNS_3 $T=5750 13320 0 0 $X=5670 $Y=13070
X56 37 M2_M1_CDNS_3 $T=6590 5910 0 0 $X=6510 $Y=5660
X57 38 M2_M1_CDNS_3 $T=7520 22860 0 0 $X=7440 $Y=22610
X58 38 M2_M1_CDNS_3 $T=7960 21030 0 0 $X=7880 $Y=20780
X59 21 M2_M1_CDNS_3 $T=8750 8160 0 0 $X=8670 $Y=7910
X60 8 M2_M1_CDNS_3 $T=8980 17010 0 0 $X=8900 $Y=16760
X61 8 M2_M1_CDNS_3 $T=10140 15570 0 0 $X=10060 $Y=15320
X62 8 M2_M1_CDNS_3 $T=10150 13320 0 0 $X=10070 $Y=13070
X63 8 M2_M1_CDNS_3 $T=10370 18740 0 0 $X=10290 $Y=18490
X64 22 M2_M1_CDNS_3 $T=10750 19470 0 0 $X=10670 $Y=19220
X65 23 M2_M1_CDNS_3 $T=11680 11800 0 0 $X=11600 $Y=11550
X66 39 M2_M1_CDNS_3 $T=12260 20780 0 0 $X=12180 $Y=20530
X67 27 M2_M1_CDNS_3 $T=13170 22790 0 0 $X=13090 $Y=22540
X68 11 M2_M1_CDNS_3 $T=13290 16990 0 0 $X=13210 $Y=16740
X69 11 M2_M1_CDNS_3 $T=14530 13310 0 0 $X=14450 $Y=13060
X70 11 M2_M1_CDNS_3 $T=14530 15600 0 0 $X=14450 $Y=15350
X71 40 M2_M1_CDNS_3 $T=14690 20780 0 0 $X=14610 $Y=20530
X72 34 M2_M1_CDNS_3 $T=15670 8330 0 0 $X=15590 $Y=8080
X73 35 M2_M1_CDNS_3 $T=16600 750 0 0 $X=16520 $Y=500
X74 23 M2_M1_CDNS_3 $T=22150 6400 0 0 $X=22070 $Y=6150
X75 26 M2_M1_CDNS_3 $T=24490 750 0 0 $X=24410 $Y=500
X76 28 M2_M1_CDNS_3 $T=26370 19410 0 0 $X=26290 $Y=19160
X77 29 M2_M1_CDNS_3 $T=26600 23000 0 0 $X=26520 $Y=22750
X78 36 M2_M1_CDNS_3 $T=28820 19250 0 0 $X=28740 $Y=19000
X79 31 M2_M1_CDNS_3 $T=29280 19170 0 0 $X=29200 $Y=18920
X80 22 M2_M1_CDNS_3 $T=33860 19960 0 90 $X=33610 $Y=19880
X81 36 M2_M1_CDNS_3 $T=34220 19150 0 0 $X=34140 $Y=18900
X82 41 M2_M1_CDNS_3 $T=35760 21100 0 0 $X=35680 $Y=20850
X83 32 M2_M1_CDNS_3 $T=35970 2380 0 0 $X=35890 $Y=2130
X84 31 M2_M1_CDNS_3 $T=39640 17490 0 0 $X=39560 $Y=17240
X85 34 M2_M1_CDNS_3 $T=43850 8260 0 0 $X=43770 $Y=8010
X86 35 M2_M1_CDNS_3 $T=43880 660 0 0 $X=43800 $Y=410
X87 36 M5_M4_CDNS_4 $T=34220 19150 0 0 $X=34140 $Y=18900
X88 29 M5_M4_CDNS_4 $T=34850 16990 0 0 $X=34770 $Y=16740
X89 36 M4_M3_CDNS_5 $T=28820 19250 0 0 $X=28740 $Y=19000
X90 36 M4_M3_CDNS_5 $T=34220 19150 0 0 $X=34140 $Y=18900
X91 1 M1_PO_CDNS_6 $T=1350 15570 0 0 $X=1250 $Y=15320
X92 1 M1_PO_CDNS_6 $T=1360 13320 0 0 $X=1260 $Y=13070
X93 7 M1_PO_CDNS_6 $T=4510 16920 0 0 $X=4410 $Y=16670
X94 7 M1_PO_CDNS_6 $T=5740 15570 0 0 $X=5640 $Y=15320
X95 7 M1_PO_CDNS_6 $T=5750 13320 0 0 $X=5650 $Y=13070
X96 37 M1_PO_CDNS_6 $T=6590 5910 0 0 $X=6490 $Y=5660
X97 38 M1_PO_CDNS_6 $T=7520 22860 0 0 $X=7420 $Y=22610
X98 38 M1_PO_CDNS_6 $T=7960 21030 0 0 $X=7860 $Y=20780
X99 8 M1_PO_CDNS_6 $T=8980 17010 0 0 $X=8880 $Y=16760
X100 8 M1_PO_CDNS_6 $T=10140 15570 0 0 $X=10040 $Y=15320
X101 8 M1_PO_CDNS_6 $T=10150 13320 0 0 $X=10050 $Y=13070
X102 8 M1_PO_CDNS_6 $T=10370 18740 0 0 $X=10270 $Y=18490
X103 22 M1_PO_CDNS_6 $T=10750 19470 0 0 $X=10650 $Y=19220
X104 39 M1_PO_CDNS_6 $T=12260 20780 0 0 $X=12160 $Y=20530
X105 11 M1_PO_CDNS_6 $T=13290 16990 0 0 $X=13190 $Y=16740
X106 11 M1_PO_CDNS_6 $T=14530 13310 0 0 $X=14430 $Y=13060
X107 11 M1_PO_CDNS_6 $T=14530 15600 0 0 $X=14430 $Y=15350
X108 40 M1_PO_CDNS_6 $T=14690 20780 0 0 $X=14590 $Y=20530
X109 34 M1_PO_CDNS_6 $T=15670 8330 0 0 $X=15570 $Y=8080
X110 35 M1_PO_CDNS_6 $T=16600 750 0 0 $X=16500 $Y=500
X111 23 M1_PO_CDNS_6 $T=22150 6400 0 0 $X=22050 $Y=6150
X112 26 M1_PO_CDNS_6 $T=24490 750 0 0 $X=24390 $Y=500
X113 31 M1_PO_CDNS_6 $T=29280 19170 0 0 $X=29180 $Y=18920
X114 36 M1_PO_CDNS_6 $T=34220 19150 0 0 $X=34120 $Y=18900
X115 41 M1_PO_CDNS_6 $T=35760 21100 0 0 $X=35660 $Y=20850
X116 32 M1_PO_CDNS_6 $T=35970 2380 0 0 $X=35870 $Y=2130
X117 1 M3_M2_CDNS_7 $T=1390 19500 0 0 $X=1310 $Y=19250
X118 19 M3_M2_CDNS_7 $T=3370 8280 0 0 $X=3290 $Y=8030
X119 20 M3_M2_CDNS_7 $T=5400 9800 0 0 $X=5320 $Y=9550
X120 7 M3_M2_CDNS_7 $T=7950 19550 0 0 $X=7870 $Y=19300
X121 24 M3_M2_CDNS_7 $T=12950 9830 0 0 $X=12870 $Y=9580
X122 25 M3_M2_CDNS_7 $T=14070 2580 0 90 $X=13820 $Y=2500
X123 26 M3_M2_CDNS_7 $T=15700 9710 0 0 $X=15620 $Y=9460
X124 11 M3_M2_CDNS_7 $T=25590 19380 0 0 $X=25510 $Y=19130
X125 27 M3_M2_CDNS_7 $T=25970 20660 0 0 $X=25890 $Y=20410
X126 30 M3_M2_CDNS_7 $T=28540 8430 0 0 $X=28460 $Y=8180
X127 30 M3_M2_CDNS_7 $T=28700 9810 0 0 $X=28620 $Y=9560
X128 33 M3_M2_CDNS_7 $T=38260 18710 0 0 $X=38180 $Y=18460
X129 32 M3_M2_CDNS_7 $T=42090 2930 0 90 $X=41840 $Y=2850
X130 2 M2_M1_CDNS_8 $T=170 4730 0 0 $X=90 $Y=4600
X131 2 M2_M1_CDNS_8 $T=180 890 0 0 $X=100 $Y=760
X132 20 M2_M1_CDNS_8 $T=4340 11800 0 0 $X=4260 $Y=11670
X133 26 M2_M1_CDNS_8 $T=8880 12210 0 0 $X=8800 $Y=12080
X134 25 M2_M1_CDNS_8 $T=13420 4530 0 0 $X=13340 $Y=4400
X135 42 M2_M1_CDNS_8 $T=17560 15460 0 0 $X=17480 $Y=15330
X136 43 M2_M1_CDNS_8 $T=21930 4780 0 0 $X=21850 $Y=4650
X137 30 M2_M1_CDNS_8 $T=29730 11900 0 0 $X=29650 $Y=11770
X138 44 M2_M1_CDNS_8 $T=31310 15530 0 0 $X=31230 $Y=15400
X139 45 M2_M1_CDNS_8 $T=35410 9580 0 0 $X=35330 $Y=9450
X140 46 M2_M1_CDNS_8 $T=41980 11840 0 0 $X=41900 $Y=11710
X141 32 M2_M1_CDNS_8 $T=43890 4790 0 0 $X=43810 $Y=4660
X142 2 M3_M2_CDNS_9 $T=160 15480 0 0 $X=80 $Y=15230
X143 2 M3_M2_CDNS_9 $T=160 21130 0 0 $X=80 $Y=20880
X144 2 M3_M2_CDNS_9 $T=170 9270 0 0 $X=90 $Y=9020
X145 2 M3_M2_CDNS_9 $T=170 13790 0 0 $X=90 $Y=13540
X146 37 M3_M2_CDNS_9 $T=500 8210 0 0 $X=420 $Y=7960
X147 1 M3_M2_CDNS_9 $T=1350 15570 0 0 $X=1270 $Y=15320
X148 1 M3_M2_CDNS_9 $T=1360 13320 0 0 $X=1280 $Y=13070
X149 39 M3_M2_CDNS_9 $T=4380 23070 0 90 $X=4130 $Y=22990
X150 19 M3_M2_CDNS_9 $T=4340 15320 0 0 $X=4260 $Y=15070
X151 47 M3_M2_CDNS_9 $T=5400 21130 0 0 $X=5320 $Y=20880
X152 7 M3_M2_CDNS_9 $T=5740 15570 0 0 $X=5660 $Y=15320
X153 7 M3_M2_CDNS_9 $T=5750 13320 0 0 $X=5670 $Y=13070
X154 37 M3_M2_CDNS_9 $T=6590 5910 0 0 $X=6510 $Y=5660
X155 38 M3_M2_CDNS_9 $T=7520 22860 0 0 $X=7440 $Y=22610
X156 38 M3_M2_CDNS_9 $T=7960 21030 0 0 $X=7880 $Y=20780
X157 48 M3_M2_CDNS_9 $T=8730 15340 0 0 $X=8650 $Y=15090
X158 8 M3_M2_CDNS_9 $T=8980 17010 0 0 $X=8900 $Y=16760
X159 8 M3_M2_CDNS_9 $T=10140 15570 0 0 $X=10060 $Y=15320
X160 8 M3_M2_CDNS_9 $T=10150 13320 0 0 $X=10070 $Y=13070
X161 24 M3_M2_CDNS_9 $T=12100 19160 0 0 $X=12020 $Y=18910
X162 39 M3_M2_CDNS_9 $T=12260 20780 0 0 $X=12180 $Y=20530
X163 49 M3_M2_CDNS_9 $T=13150 15340 0 0 $X=13070 $Y=15090
X164 40 M3_M2_CDNS_9 $T=14690 20780 0 0 $X=14610 $Y=20530
X165 34 M3_M2_CDNS_9 $T=15670 8330 0 0 $X=15590 $Y=8080
X166 35 M3_M2_CDNS_9 $T=16600 750 0 0 $X=16520 $Y=500
X167 40 M3_M2_CDNS_9 $T=17570 22850 0 0 $X=17490 $Y=22600
X168 36 M3_M2_CDNS_9 $T=22230 22840 0 0 $X=22150 $Y=22590
X169 36 M3_M2_CDNS_9 $T=28820 20830 0 0 $X=28740 $Y=20580
X170 41 M3_M2_CDNS_9 $T=35370 22940 0 0 $X=35290 $Y=22690
X171 19 M3_M2_CDNS_10 $T=4340 13390 0 0 $X=4260 $Y=13260
X172 47 M3_M2_CDNS_10 $T=7370 12440 0 0 $X=7290 $Y=12310
X173 47 M3_M2_CDNS_10 $T=8600 9080 0 0 $X=8520 $Y=8950
X174 8 M3_M2_CDNS_10 $T=10370 18740 0 0 $X=10290 $Y=18610
X175 24 M3_M2_CDNS_10 $T=13190 12020 0 0 $X=13110 $Y=11890
X176 43 M3_M2_CDNS_10 $T=19690 2880 0 90 $X=19560 $Y=2800
X177 27 M3_M2_CDNS_10 $T=26840 17540 0 90 $X=26710 $Y=17460
X178 41 M3_M2_CDNS_10 $T=35760 21100 0 0 $X=35680 $Y=20970
X179 29 M4_M3_CDNS_11 $T=34850 16990 0 0 $X=34770 $Y=16740
X180 1 M4_M3_CDNS_12 $T=1390 21140 0 0 $X=1310 $Y=21010
X181 19 M4_M3_CDNS_12 $T=3650 6110 0 0 $X=3570 $Y=5980
X182 20 M4_M3_CDNS_12 $T=6680 2460 0 0 $X=6600 $Y=2330
X183 27 M4_M3_CDNS_12 $T=13170 22790 0 0 $X=13090 $Y=22660
X184 24 M4_M3_CDNS_12 $T=13680 4950 0 0 $X=13600 $Y=4820
X185 11 M4_M3_CDNS_12 $T=14530 13310 0 0 $X=14450 $Y=13180
X186 11 M4_M3_CDNS_12 $T=14530 15600 0 0 $X=14450 $Y=15470
X187 25 M4_M3_CDNS_12 $T=21870 1570 0 0 $X=21790 $Y=1440
X188 21 M4_M3_CDNS_12 $T=23120 3950 0 0 $X=23040 $Y=3820
X189 28 M4_M3_CDNS_12 $T=28320 12210 0 0 $X=28240 $Y=12080
X190 35 M4_M3_CDNS_12 $T=28540 230 0 90 $X=28410 $Y=150
X191 34 M4_M3_CDNS_12 $T=28550 7610 0 90 $X=28420 $Y=7530
X192 22 M4_M3_CDNS_12 $T=33860 19960 0 90 $X=33730 $Y=19880
X193 2 M2_M1_CDNS_13 $T=160 15480 0 0 $X=80 $Y=15230
X194 2 M2_M1_CDNS_13 $T=160 21130 0 0 $X=80 $Y=20880
X195 2 M2_M1_CDNS_13 $T=170 9270 0 0 $X=90 $Y=9020
X196 2 M2_M1_CDNS_13 $T=170 13790 0 0 $X=90 $Y=13540
X197 37 M2_M1_CDNS_13 $T=500 8210 0 0 $X=420 $Y=7960
X198 39 M2_M1_CDNS_13 $T=4380 23070 0 90 $X=4130 $Y=22990
X199 19 M2_M1_CDNS_13 $T=4340 15320 0 0 $X=4260 $Y=15070
X200 47 M2_M1_CDNS_13 $T=5400 21130 0 0 $X=5320 $Y=20880
X201 48 M2_M1_CDNS_13 $T=8730 15340 0 0 $X=8650 $Y=15090
X202 24 M2_M1_CDNS_13 $T=12100 19160 0 0 $X=12020 $Y=18910
X203 49 M2_M1_CDNS_13 $T=13150 15340 0 0 $X=13070 $Y=15090
X204 40 M2_M1_CDNS_13 $T=17570 22850 0 0 $X=17490 $Y=22600
X205 36 M2_M1_CDNS_13 $T=22230 22840 0 0 $X=22150 $Y=22590
X206 36 M2_M1_CDNS_13 $T=28820 20830 0 0 $X=28740 $Y=20580
X207 41 M2_M1_CDNS_13 $T=35370 22940 0 0 $X=35290 $Y=22690
X208 33 M2_M1_CDNS_13 $T=46340 18970 0 0 $X=46260 $Y=18720
X209 36 M5_M4_CDNS_14 $T=28820 19250 0 0 $X=28740 $Y=19120
X210 29 M5_M4_CDNS_14 $T=35550 19590 0 0 $X=35470 $Y=19460
X211 1 M1_PO_CDNS_15 $T=1390 17230 0 0 $X=1290 $Y=16980
X212 1 M1_PO_CDNS_15 $T=1390 24660 0 0 $X=1290 $Y=24410
X213 3 M1_PO_CDNS_15 $T=2770 22320 0 90 $X=2520 $Y=22220
X214 5 M1_PO_CDNS_15 $T=2650 13610 0 0 $X=2550 $Y=13360
X215 4 M1_PO_CDNS_15 $T=2750 17050 0 0 $X=2650 $Y=16800
X216 1 M1_PO_CDNS_15 $T=4410 23850 0 0 $X=4310 $Y=23600
X217 4 M1_PO_CDNS_15 $T=5790 16970 0 0 $X=5690 $Y=16720
X218 9 M1_PO_CDNS_15 $T=7290 23970 0 90 $X=7040 $Y=23870
X219 5 M1_PO_CDNS_15 $T=7180 13450 0 0 $X=7080 $Y=13200
X220 3 M1_PO_CDNS_15 $T=8720 22330 0 90 $X=8470 $Y=22230
X221 3 M1_PO_CDNS_15 $T=9910 24890 0 90 $X=9660 $Y=24790
X222 4 M1_PO_CDNS_15 $T=10210 17010 0 0 $X=10110 $Y=16760
X223 7 M1_PO_CDNS_15 $T=11550 22710 0 0 $X=11450 $Y=22460
X224 5 M1_PO_CDNS_15 $T=11730 13390 0 0 $X=11630 $Y=13140
X225 9 M1_PO_CDNS_15 $T=13230 23970 0 90 $X=12980 $Y=23870
X226 4 M1_PO_CDNS_15 $T=14630 17040 0 0 $X=14530 $Y=16790
X227 7 M1_PO_CDNS_15 $T=15790 22330 0 90 $X=15540 $Y=22230
X228 5 M1_PO_CDNS_15 $T=15980 13520 0 0 $X=15880 $Y=13270
X229 3 M1_PO_CDNS_15 $T=17780 24480 0 0 $X=17680 $Y=24230
X230 8 M1_PO_CDNS_15 $T=20560 22320 0 90 $X=20310 $Y=22220
X231 9 M1_PO_CDNS_15 $T=22240 23950 0 0 $X=22140 $Y=23700
X232 8 M1_PO_CDNS_15 $T=24880 22320 0 90 $X=24630 $Y=22220
X233 3 M1_PO_CDNS_15 $T=26710 24400 0 0 $X=26610 $Y=24150
X234 30 M1_PO_CDNS_15 $T=28540 6330 0 0 $X=28440 $Y=6080
X235 11 M1_PO_CDNS_15 $T=29350 22530 0 0 $X=29250 $Y=22280
X236 42 M1_PO_CDNS_15 $T=29800 13490 0 0 $X=29700 $Y=13240
X237 9 M1_PO_CDNS_15 $T=31140 23850 0 0 $X=31040 $Y=23600
X238 44 M1_PO_CDNS_15 $T=31170 13680 0 0 $X=31070 $Y=13430
X239 33 M1_PO_CDNS_15 $T=31860 16950 0 0 $X=31760 $Y=16700
X240 11 M1_PO_CDNS_15 $T=33650 22300 0 90 $X=33400 $Y=22200
X241 46 M1_PO_CDNS_15 $T=35890 9730 0 0 $X=35790 $Y=9480
X242 1 M2_M1_CDNS_17 $T=1390 17230 0 0 $X=1310 $Y=16980
X243 1 M2_M1_CDNS_17 $T=1390 24660 0 0 $X=1310 $Y=24410
X244 3 M2_M1_CDNS_17 $T=2770 22320 0 90 $X=2520 $Y=22240
X245 5 M2_M1_CDNS_17 $T=2650 13610 0 0 $X=2570 $Y=13360
X246 4 M2_M1_CDNS_17 $T=2750 17050 0 0 $X=2670 $Y=16800
X247 1 M2_M1_CDNS_17 $T=4410 23850 0 0 $X=4330 $Y=23600
X248 4 M2_M1_CDNS_17 $T=5790 16970 0 0 $X=5710 $Y=16720
X249 9 M2_M1_CDNS_17 $T=7290 23970 0 90 $X=7040 $Y=23890
X250 5 M2_M1_CDNS_17 $T=7180 13450 0 0 $X=7100 $Y=13200
X251 3 M2_M1_CDNS_17 $T=8720 22330 0 90 $X=8470 $Y=22250
X252 3 M2_M1_CDNS_17 $T=9910 24890 0 90 $X=9660 $Y=24810
X253 4 M2_M1_CDNS_17 $T=10210 17010 0 0 $X=10130 $Y=16760
X254 7 M2_M1_CDNS_17 $T=11550 22710 0 0 $X=11470 $Y=22460
X255 5 M2_M1_CDNS_17 $T=11730 13390 0 0 $X=11650 $Y=13140
X256 9 M2_M1_CDNS_17 $T=13230 23970 0 90 $X=12980 $Y=23890
X257 4 M2_M1_CDNS_17 $T=14630 17040 0 0 $X=14550 $Y=16790
X258 7 M2_M1_CDNS_17 $T=15790 22330 0 90 $X=15540 $Y=22250
X259 5 M2_M1_CDNS_17 $T=15980 13520 0 0 $X=15900 $Y=13270
X260 3 M2_M1_CDNS_17 $T=17780 24480 0 0 $X=17700 $Y=24230
X261 8 M2_M1_CDNS_17 $T=20560 22320 0 90 $X=20310 $Y=22240
X262 9 M2_M1_CDNS_17 $T=22240 23950 0 0 $X=22160 $Y=23700
X263 8 M2_M1_CDNS_17 $T=24880 22320 0 90 $X=24630 $Y=22240
X264 3 M2_M1_CDNS_17 $T=26710 24400 0 0 $X=26630 $Y=24150
X265 30 M2_M1_CDNS_17 $T=28540 6330 0 0 $X=28460 $Y=6080
X266 11 M2_M1_CDNS_17 $T=29350 22530 0 0 $X=29270 $Y=22280
X267 42 M2_M1_CDNS_17 $T=29800 13490 0 0 $X=29720 $Y=13240
X268 9 M2_M1_CDNS_17 $T=31140 23850 0 0 $X=31060 $Y=23600
X269 44 M2_M1_CDNS_17 $T=31170 13680 0 0 $X=31090 $Y=13430
X270 33 M2_M1_CDNS_17 $T=31860 16950 0 0 $X=31780 $Y=16700
X271 11 M2_M1_CDNS_17 $T=33650 22300 0 90 $X=33400 $Y=22220
X272 46 M2_M1_CDNS_17 $T=35890 9730 0 0 $X=35810 $Y=9480
X273 1 6 2 5 20 77 AND $T=40 14460 1 0 $X=50 $Y=10660
X274 1 6 2 4 19 76 AND $T=40 14420 0 0 $X=50 $Y=14420
X275 1 6 2 3 39 75 AND $T=40 21740 0 0 $X=50 $Y=21740
X276 7 6 2 5 26 80 AND $T=4440 14460 1 0 $X=4450 $Y=10660
X277 7 6 2 4 48 79 AND $T=4440 14420 0 0 $X=4450 $Y=14420
X278 1 6 2 9 38 78 AND $T=4440 21740 0 0 $X=4450 $Y=21740
X279 8 6 2 5 23 83 AND $T=8840 14460 1 0 $X=8850 $Y=10660
X280 8 6 2 4 49 82 AND $T=8840 14420 0 0 $X=8850 $Y=14420
X281 3 6 2 7 27 81 AND $T=8840 21740 0 0 $X=8850 $Y=21740
X282 11 6 2 5 50 93 AND $T=13240 14460 1 0 $X=13250 $Y=10660
X283 11 6 2 4 42 92 AND $T=13240 14420 0 0 $X=13250 $Y=14420
X284 9 6 2 7 40 91 AND $T=13240 21740 0 0 $X=13250 $Y=21740
X285 3 6 2 8 36 104 AND $T=17880 21740 0 0 $X=17890 $Y=21740
X286 9 6 2 8 29 126 AND $T=22280 21740 0 0 $X=22290 $Y=21740
X287 3 6 2 11 14 127 AND $T=26680 21740 0 0 $X=26690 $Y=21740
X288 9 6 2 11 41 131 AND $T=31080 21740 0 0 $X=31090 $Y=21740
X289 38 2 6 22 47 24 73 74 225 half_adder $T=50 21780 1 0 $X=50 $Y=17980
X290 50 2 6 45 13 30 102 103 228 half_adder $T=17640 14460 1 0 $X=17640 $Y=10660
X291 42 2 6 44 17 46 129 130 237 half_adder $T=29830 14460 1 0 $X=29830 $Y=10660
X292 36 2 6 41 18 33 133 134 238 half_adder $T=34210 21780 1 0 $X=34210 $Y=17980
X293 47 6 48 2 34 21 37 67 70 71
+ 65 66 68 69 223 224 full_adder1_small $T=22270 7090 1 180 $X=20 $Y=7100
X294 20 6 43 2 35 10 12 60 63 64
+ 58 59 61 62 221 222 full_adder1_small $T=30 -230 0 0 $X=50 $Y=-220
X295 19 6 24 2 37 25 43 53 56 57
+ 51 52 54 55 219 220 full_adder1_small $T=30 7150 1 0 $X=50 $Y=3340
X296 39 6 40 2 31 28 22 86 89 90
+ 84 85 87 88 226 227 full_adder1_small $T=12230 21790 1 0 $X=12250 $Y=17980
X297 29 6 27 2 33 44 31 96 99 100
+ 94 95 97 98 229 230 full_adder1_small $T=17850 14410 0 0 $X=17870 $Y=14420
X298 26 6 25 2 32 15 35 121 124 125
+ 119 120 122 123 235 236 full_adder1_small $T=21990 -230 0 0 $X=22010 $Y=-220
X299 23 6 21 2 30 16 32 114 117 118
+ 112 113 115 116 233 234 full_adder1_small $T=21990 7150 1 0 $X=22010 $Y=3340
X300 49 6 28 2 46 45 34 107 110 111
+ 105 106 108 109 231 232 full_adder1_small $T=21990 7090 0 0 $X=22010 $Y=7100
M0 77 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=11610 $dt=1
M1 76 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=16790 $dt=1
M2 75 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=24110 $dt=1
M3 73 38 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=16.2188 scb=0.0173423 scc=0.000698846 $X=750 $Y=18640 $dt=1
M4 58 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=2120 $dt=1
M5 51 19 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=4320 $dt=1
M6 37 71 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=1070 $Y=9450 $dt=1
M7 6 70 37 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=1480 $Y=9450 $dt=1
M8 59 43 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=2120 $dt=1
M9 52 24 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=4320 $dt=1
M10 77 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=11600 $dt=1
M11 76 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=16800 $dt=1
M12 75 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=24120 $dt=1
M13 221 43 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=1880 $dt=1
M14 219 24 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=4080 $dt=1
M15 20 77 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=11580 $dt=1
M16 19 76 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=16820 $dt=1
M17 39 75 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=24140 $dt=1
M18 71 48 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=3910 $Y=9450 $dt=1
M19 60 58 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=1940 $dt=1
M20 53 51 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=4020 $dt=1
M21 6 47 71 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=4320 $Y=9450 $dt=1
M22 60 59 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=1940 $dt=1
M23 53 52 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=4020 $dt=1
M24 80 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=11610 $dt=1
M25 79 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=16790 $dt=1
M26 78 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=24110 $dt=1
M27 221 20 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=1940 $dt=1
M28 219 19 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=4020 $dt=1
M29 47 22 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=6190 $Y=18700 $dt=1
M30 80 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=11600 $dt=1
M31 79 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=16800 $dt=1
M32 78 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=24120 $dt=1
M33 70 67 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=6890 $Y=9230 $dt=1
M34 6 34 70 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=7300 $Y=9230 $dt=1
M35 47 38 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=7300 $Y=18660 $dt=1
M36 61 35 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=2120 $dt=1
M37 54 37 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=4320 $dt=1
M38 26 80 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=11580 $dt=1
M39 48 79 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=16820 $dt=1
M40 38 78 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=24140 $dt=1
M41 74 38 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=8540 $Y=18930 $dt=1
M42 62 60 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=2120 $dt=1
M43 55 53 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=4320 $dt=1
M44 6 34 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=9370 $Y=9260 $dt=1
M45 83 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=11610 $dt=1
M46 82 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=16790 $dt=1
M47 81 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=24110 $dt=1
M48 74 22 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=9780 $Y=18920 $dt=1
M49 222 60 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=1880 $dt=1
M50 220 53 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=4080 $dt=1
M51 224 69 21 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10330 $Y=9260 $dt=1
M52 83 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=11600 $dt=1
M53 82 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=16800 $dt=1
M54 81 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=24120 $dt=1
M55 10 61 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=1940 $dt=1
M56 25 54 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=4020 $dt=1
M57 224 68 21 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11290 $Y=9260 $dt=1
M58 24 74 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=11460 $Y=18900 $dt=1
M59 10 62 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=1940 $dt=1
M60 25 55 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=4020 $dt=1
M61 6 67 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=12260 $Y=9200 $dt=1
M62 23 83 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=11580 $dt=1
M63 49 82 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=16820 $dt=1
M64 27 81 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=24140 $dt=1
M65 222 35 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=1940 $dt=1
M66 220 37 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=4020 $dt=1
M67 84 39 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13020 $Y=18960 $dt=1
M68 6 67 69 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13590 $Y=9440 $dt=1
M69 93 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=11610 $dt=1
M70 92 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=16790 $dt=1
M71 91 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=24110 $dt=1
M72 85 40 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13980 $Y=18960 $dt=1
M73 6 34 68 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=14550 $Y=9440 $dt=1
M74 63 35 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=1910 $dt=1
M75 56 37 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=4050 $dt=1
M76 93 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=11600 $dt=1
M77 92 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=16800 $dt=1
M78 91 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=24120 $dt=1
M79 226 40 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=15310 $Y=18720 $dt=1
M80 6 60 63 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=1910 $dt=1
M81 6 53 56 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=4050 $dt=1
M82 6 47 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16210 $Y=9260 $dt=1
M83 86 84 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16280 $Y=18660 $dt=1
M84 50 93 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=11580 $dt=1
M85 42 92 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=16820 $dt=1
M86 40 91 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=24140 $dt=1
M87 223 66 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17170 $Y=9260 $dt=1
M88 86 85 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17240 $Y=18660 $dt=1
M89 64 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=2130 $dt=1
M90 57 19 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=4310 $dt=1
M91 223 65 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18130 $Y=9260 $dt=1
M92 226 39 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18200 $Y=18660 $dt=1
M93 6 43 64 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=2130 $dt=1
M94 6 24 57 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=4310 $dt=1
M95 102 50 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=18340 $Y=11320 $dt=1
M96 104 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=18580 $Y=24110 $dt=1
M97 94 29 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=18640 $Y=16760 $dt=1
M98 6 48 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=19100 $Y=9200 $dt=1
M99 95 27 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19600 $Y=16760 $dt=1
M100 104 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=19820 $Y=24120 $dt=1
M101 87 31 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19860 $Y=18960 $dt=1
M102 6 48 66 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20430 $Y=9440 $dt=1
M103 12 63 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=2130 $dt=1
M104 43 56 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=4310 $dt=1
M105 88 86 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20820 $Y=18960 $dt=1
M106 229 27 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=20930 $Y=16520 $dt=1
M107 6 64 12 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=2130 $dt=1
M108 6 57 43 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=4310 $dt=1
M109 6 47 65 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=21390 $Y=9440 $dt=1
M110 36 104 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=21500 $Y=24140 $dt=1
M111 96 94 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=21900 $Y=16580 $dt=1
M112 227 86 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=22150 $Y=18720 $dt=1
M113 119 26 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=2120 $dt=1
M114 112 23 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=4320 $dt=1
M115 105 49 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=9440 $dt=1
M116 96 95 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=22860 $Y=16580 $dt=1
M117 126 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=22980 $Y=24110 $dt=1
M118 28 87 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23120 $Y=18660 $dt=1
M119 120 25 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=2120 $dt=1
M120 113 21 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=4320 $dt=1
M121 106 28 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=9440 $dt=1
M122 13 45 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=23780 $Y=11380 $dt=1
M123 229 29 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23820 $Y=16580 $dt=1
M124 28 88 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24080 $Y=18660 $dt=1
M125 126 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=24220 $Y=24120 $dt=1
M126 13 50 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24890 $Y=11340 $dt=1
M127 227 31 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=25040 $Y=18660 $dt=1
M128 235 25 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=1880 $dt=1
M129 233 21 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=4080 $dt=1
M130 231 28 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=9200 $dt=1
M131 97 33 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=25480 $Y=16760 $dt=1
M132 29 126 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=25900 $Y=24140 $dt=1
M133 121 119 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=1940 $dt=1
M134 114 112 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=4020 $dt=1
M135 107 105 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=9260 $dt=1
M136 103 50 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26130 $Y=11610 $dt=1
M137 98 96 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=26440 $Y=16760 $dt=1
M138 121 120 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=1940 $dt=1
M139 114 113 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=4020 $dt=1
M140 107 106 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=9260 $dt=1
M141 89 31 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27110 $Y=18690 $dt=1
M142 103 45 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27370 $Y=11600 $dt=1
M143 127 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=27380 $Y=24110 $dt=1
M144 6 86 89 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27520 $Y=18690 $dt=1
M145 230 96 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=27770 $Y=16520 $dt=1
M146 235 26 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=1940 $dt=1
M147 233 23 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=4020 $dt=1
M148 231 49 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=9260 $dt=1
M149 127 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=28620 $Y=24120 $dt=1
M150 44 97 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28740 $Y=16580 $dt=1
M151 30 103 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=29050 $Y=11580 $dt=1
M152 122 32 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=2120 $dt=1
M153 115 30 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=4320 $dt=1
M154 108 46 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=9440 $dt=1
M155 44 98 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=29700 $Y=16580 $dt=1
M156 90 39 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30090 $Y=18950 $dt=1
M157 14 127 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=30300 $Y=24140 $dt=1
M158 6 40 90 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30500 $Y=18950 $dt=1
M159 129 42 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=30530 $Y=11320 $dt=1
M160 123 121 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=2120 $dt=1
M161 116 114 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=4320 $dt=1
M162 109 107 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=9440 $dt=1
M163 230 33 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=30660 $Y=16580 $dt=1
M164 131 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=31780 $Y=24110 $dt=1
M165 236 121 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=1880 $dt=1
M166 234 114 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=4080 $dt=1
M167 232 107 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=9200 $dt=1
M168 99 33 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=32730 $Y=16550 $dt=1
M169 15 122 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=1940 $dt=1
M170 16 115 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=4020 $dt=1
M171 45 108 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=9260 $dt=1
M172 22 89 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=32930 $Y=18950 $dt=1
M173 131 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=33020 $Y=24120 $dt=1
M174 6 96 99 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=33140 $Y=16550 $dt=1
M175 6 90 22 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=33340 $Y=18950 $dt=1
M176 15 123 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=1940 $dt=1
M177 16 116 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=4020 $dt=1
M178 45 109 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=9260 $dt=1
M179 41 131 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=34700 $Y=24140 $dt=1
M180 236 32 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=1940 $dt=1
M181 234 30 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=4020 $dt=1
M182 232 46 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=9260 $dt=1
M183 133 36 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=34910 $Y=18640 $dt=1
M184 100 29 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=35710 $Y=16770 $dt=1
M185 17 44 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=35970 $Y=11380 $dt=1
M186 6 27 100 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=36120 $Y=16770 $dt=1
M187 124 32 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=1910 $dt=1
M188 117 30 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=4050 $dt=1
M189 110 46 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=9230 $dt=1
M190 17 42 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=37080 $Y=11340 $dt=1
M191 6 121 124 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=1910 $dt=1
M192 6 114 117 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=4050 $dt=1
M193 6 107 110 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=9230 $dt=1
M194 130 42 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=38320 $Y=11610 $dt=1
M195 31 99 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=38550 $Y=16770 $dt=1
M196 6 100 31 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=38960 $Y=16770 $dt=1
M197 130 44 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=39560 $Y=11600 $dt=1
M198 125 26 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=2130 $dt=1
M199 118 23 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=4310 $dt=1
M200 111 49 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=9450 $dt=1
M201 6 25 125 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=2130 $dt=1
M202 6 21 118 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=4310 $dt=1
M203 6 28 111 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=9450 $dt=1
M204 18 41 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.2705 scb=0.0126902 scc=0.000796523 $X=40350 $Y=18700 $dt=1
M205 46 130 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=41240 $Y=11580 $dt=1
M206 18 36 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=41460 $Y=18660 $dt=1
M207 35 124 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=2130 $dt=1
M208 32 117 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=4310 $dt=1
M209 34 110 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=42690 $Y=9450 $dt=1
M210 134 36 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42700 $Y=18930 $dt=1
M211 6 125 35 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=2130 $dt=1
M212 6 118 32 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=4310 $dt=1
M213 6 111 34 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=43100 $Y=9450 $dt=1
M214 134 41 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43940 $Y=18920 $dt=1
M215 33 134 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=45620 $Y=18900 $dt=1
.ends multiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_31                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_31 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_31

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_32                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_32 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_32

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_43                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_43 1 2 3 5 6 8
*.DEVICECLIMB
** N=14 EP=6 FDC=2
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=810 $Y=710 $dt=0
M1 8 6 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=4640 $Y=580 $dt=0
.ends cellTmpl_CDNS_43

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_44                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_44 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_44

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_45                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_45 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_45

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=12
X0 7 M2_M1_CDNS_3 $T=250 -3000 0 0 $X=170 $Y=-3250
X1 7 M2_M1_CDNS_3 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X2 7 M1_PO_CDNS_6 $T=250 -3000 0 0 $X=150 $Y=-3250
X3 7 M1_PO_CDNS_6 $T=2620 -2730 0 0 $X=2520 $Y=-2980
X4 7 M3_M2_CDNS_9 $T=250 -3000 0 0 $X=170 $Y=-3250
X5 7 M3_M2_CDNS_9 $T=960 -2040 0 0 $X=880 $Y=-2290
X6 7 M3_M2_CDNS_9 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X7 7 M2_M1_CDNS_13 $T=960 -2040 0 0 $X=880 $Y=-2290
X8 1 M1_PO_CDNS_15 $T=1300 -3500 0 0 $X=1200 $Y=-3750
X9 1 M1_PO_CDNS_15 $T=2660 -4240 0 0 $X=2560 $Y=-4490
X10 1 M1_PO_CDNS_16 $T=680 -3550 0 0 $X=580 $Y=-3670
X11 2 M1_PO_CDNS_16 $T=1300 -2090 0 0 $X=1200 $Y=-2210
X12 5 M1_PO_CDNS_16 $T=4040 -3180 0 0 $X=3940 $Y=-3300
X13 8 M1_PO_CDNS_16 $T=4300 -3670 0 90 $X=4180 $Y=-3770
X14 1 M2_M1_CDNS_17 $T=1300 -3500 0 0 $X=1220 $Y=-3750
X15 1 M2_M1_CDNS_17 $T=2660 -4240 0 0 $X=2580 $Y=-4490
X16 4 7 9 4 nmos1v_CDNS_31 $T=1990 -4420 0 0 $X=1790 $Y=-4620
X17 8 5 10 4 nmos1v_CDNS_31 $T=3370 -4430 0 0 $X=3170 $Y=-4630
X18 8 2 9 4 nmos1v_CDNS_32 $T=1780 -4420 0 0 $X=1360 $Y=-4620
X19 4 1 10 4 nmos1v_CDNS_32 $T=3160 -4430 0 0 $X=2740 $Y=-4630
X20 3 4 1 7 8 6 cellTmpl_CDNS_43 $T=-60 -5080 0 0 $X=-180 $Y=-5220
X21 3 1 11 4 3 pmos1v_CDNS_44 $T=1990 -3120 0 0 $X=1790 $Y=-3320
X22 8 5 12 4 3 pmos1v_CDNS_44 $T=3370 -3190 0 0 $X=3170 $Y=-3390
X23 8 2 11 4 3 pmos1v_CDNS_45 $T=1780 -3120 0 0 $X=1360 $Y=-3320
X24 3 7 12 4 3 pmos1v_CDNS_45 $T=3160 -3190 0 0 $X=2740 $Y=-3390
M0 9 2 8 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1780 $Y=-4420 $dt=0
M1 4 7 9 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1990 $Y=-4420 $dt=0
M2 10 1 4 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3160 $Y=-4430 $dt=0
M3 8 5 10 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3370 $Y=-4430 $dt=0
M4 7 1 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=750 $Y=-2850 $dt=1
M5 11 2 8 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1780 $Y=-3120 $dt=1
M6 3 1 11 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1990 $Y=-3120 $dt=1
M7 12 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3160 $Y=-3190 $dt=1
M8 8 5 12 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3370 $Y=-3190 $dt=1
M9 6 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.2373 scb=0.0194294 scc=0.00149528 $X=4580 $Y=-3180 $dt=1
.ends MUX_2to1___2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FA_4bit                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FA_4bit 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19
** N=83 EP=19 FDC=144
X0 17 M4_M3_CDNS_1 $T=14030 6120 0 0 $X=13950 $Y=5870
X1 18 M4_M3_CDNS_1 $T=16960 11880 0 0 $X=16880 $Y=11630
X2 17 M4_M3_CDNS_1 $T=19730 4760 0 0 $X=19650 $Y=4510
X3 18 M4_M3_CDNS_1 $T=22610 11350 0 0 $X=22530 $Y=11100
X4 17 M3_M2_CDNS_2 $T=14030 6120 0 0 $X=13950 $Y=5870
X5 18 M3_M2_CDNS_2 $T=16960 11880 0 0 $X=16880 $Y=11630
X6 18 M3_M2_CDNS_2 $T=22610 11350 0 0 $X=22530 $Y=11100
X7 17 M2_M1_CDNS_3 $T=14030 6120 0 0 $X=13950 $Y=5870
X8 18 M2_M1_CDNS_3 $T=16960 11880 0 0 $X=16880 $Y=11630
X9 19 M2_M1_CDNS_3 $T=18840 8310 0 0 $X=18760 $Y=8060
X10 18 M2_M1_CDNS_3 $T=22610 11350 0 0 $X=22530 $Y=11100
X11 17 M1_PO_CDNS_6 $T=14030 6120 0 0 $X=13930 $Y=5870
X12 18 M1_PO_CDNS_6 $T=16960 11880 0 0 $X=16860 $Y=11630
X13 19 M1_PO_CDNS_6 $T=18840 8310 0 0 $X=18740 $Y=8060
X14 17 M3_M2_CDNS_7 $T=19730 4760 0 0 $X=19650 $Y=4510
X15 5 M2_M1_CDNS_8 $T=-80 3540 0 0 $X=-160 $Y=3410
X16 5 M2_M1_CDNS_8 $T=-80 10890 0 0 $X=-160 $Y=10760
X17 17 M2_M1_CDNS_8 $T=21770 2020 0 0 $X=21690 $Y=1890
X18 19 M2_M1_CDNS_8 $T=21770 5100 0 0 $X=21690 $Y=4970
X19 19 M3_M2_CDNS_9 $T=18840 8310 0 0 $X=18760 $Y=8060
X20 19 M3_M2_CDNS_10 $T=21980 9220 0 0 $X=21900 $Y=9090
X21 6 5 1 7 11 12 17 43 46 47
+ 41 42 44 45 82 83 full_adder1_small $T=-90 -130 0 0 $X=-70 $Y=-120
X22 8 5 2 7 17 13 19 36 39 40
+ 34 35 37 38 80 81 full_adder1_small $T=-90 7250 1 0 $X=-70 $Y=3440
X23 9 5 3 7 19 14 18 29 32 33
+ 27 28 30 31 78 79 full_adder1_small $T=-90 7190 0 0 $X=-70 $Y=7200
X24 10 5 4 7 18 15 16 22 25 26
+ 20 21 23 24 76 77 full_adder1_small $T=-90 14570 1 0 $X=-70 $Y=10760
M0 41 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=2220 $dt=1
M1 34 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=4420 $dt=1
M2 27 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=9540 $dt=1
M3 20 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=11740 $dt=1
M4 42 1 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=2220 $dt=1
M5 35 2 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=4420 $dt=1
M6 28 3 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=9540 $dt=1
M7 21 4 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=11740 $dt=1
M8 82 1 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=1980 $dt=1
M9 80 2 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=4180 $dt=1
M10 78 3 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=9300 $dt=1
M11 76 4 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=11500 $dt=1
M12 43 41 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=2040 $dt=1
M13 36 34 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=4120 $dt=1
M14 29 27 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=9360 $dt=1
M15 22 20 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=11440 $dt=1
M16 43 42 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=2040 $dt=1
M17 36 35 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=4120 $dt=1
M18 29 28 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=9360 $dt=1
M19 22 21 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=11440 $dt=1
M20 82 6 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=2040 $dt=1
M21 80 8 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=4120 $dt=1
M22 78 9 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=9360 $dt=1
M23 76 10 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=11440 $dt=1
M24 44 11 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=2220 $dt=1
M25 37 17 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=4420 $dt=1
M26 30 19 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=9540 $dt=1
M27 23 18 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=11740 $dt=1
M28 45 43 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=2220 $dt=1
M29 38 36 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=4420 $dt=1
M30 31 29 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=9540 $dt=1
M31 24 22 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=11740 $dt=1
M32 83 43 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=1980 $dt=1
M33 81 36 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=4180 $dt=1
M34 79 29 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=9300 $dt=1
M35 77 22 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=11500 $dt=1
M36 12 44 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=2040 $dt=1
M37 13 37 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=4120 $dt=1
M38 14 30 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=9360 $dt=1
M39 15 23 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=11440 $dt=1
M40 12 45 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=2040 $dt=1
M41 13 38 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=4120 $dt=1
M42 14 31 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=9360 $dt=1
M43 15 24 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=11440 $dt=1
M44 83 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=2040 $dt=1
M45 81 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=4120 $dt=1
M46 79 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=9360 $dt=1
M47 77 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=11440 $dt=1
M48 46 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=2010 $dt=1
M49 39 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=4150 $dt=1
M50 32 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=9330 $dt=1
M51 25 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=11470 $dt=1
M52 5 43 46 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=2010 $dt=1
M53 5 36 39 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=4150 $dt=1
M54 5 29 32 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=9330 $dt=1
M55 5 22 25 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=11470 $dt=1
M56 47 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=2230 $dt=1
M57 40 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=4410 $dt=1
M58 33 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=9550 $dt=1
M59 26 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=11730 $dt=1
M60 5 1 47 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=2230 $dt=1
M61 5 2 40 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=4410 $dt=1
M62 5 3 33 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=9550 $dt=1
M63 5 4 26 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=11730 $dt=1
M64 17 46 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=2230 $dt=1
M65 19 39 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=4410 $dt=1
M66 18 32 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=9550 $dt=1
M67 16 25 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=11730 $dt=1
M68 5 47 17 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=2230 $dt=1
M69 5 40 19 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=4410 $dt=1
M70 5 33 18 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=9550 $dt=1
M71 5 26 16 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=11730 $dt=1
.ends FA_4bit

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small 1 2 3 4
** N=4 EP=4 FDC=2
X0 1 M1_PO_CDNS_16 $T=950 1780 0 90 $X=830 $Y=1680
X1 2 3 cellTmpl_CDNS_18 $T=120 140 0 0 $X=0 $Y=0
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7353 scb=0.0117274 scc=0.000445561 $X=1070 $Y=980 $dt=0
M1 4 1 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8675 scb=0.0146094 scc=0.000688105 $X=1070 $Y=2220 $dt=1
.ends INV_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 10badder                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 10badder 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59
** N=267 EP=59 FDC=516
X0 35 M4_M3_CDNS_1 $T=51080 34160 0 0 $X=51000 $Y=33910
X1 36 M4_M3_CDNS_1 $T=56340 32800 0 0 $X=56260 $Y=32550
X2 37 M4_M3_CDNS_1 $T=56340 47440 0 0 $X=56260 $Y=47190
X3 38 M4_M3_CDNS_1 $T=57240 50840 0 0 $X=57160 $Y=50590
X4 39 M4_M3_CDNS_1 $T=72650 52420 0 90 $X=72400 $Y=52340
X5 35 M4_M3_CDNS_1 $T=78550 36430 0 0 $X=78470 $Y=36180
X6 39 M4_M3_CDNS_1 $T=79400 52420 0 90 $X=79150 $Y=52340
X7 36 M4_M3_CDNS_1 $T=86760 34460 0 0 $X=86680 $Y=34210
X8 37 M4_M3_CDNS_1 $T=86760 49100 0 0 $X=86680 $Y=48850
X9 35 M3_M2_CDNS_2 $T=51080 34160 0 0 $X=51000 $Y=33910
X10 36 M3_M2_CDNS_2 $T=56340 32800 0 0 $X=56260 $Y=32550
X11 37 M3_M2_CDNS_2 $T=56340 47440 0 0 $X=56260 $Y=47190
X12 38 M3_M2_CDNS_2 $T=57240 50840 0 0 $X=57160 $Y=50590
X13 39 M3_M2_CDNS_2 $T=72650 52420 0 90 $X=72400 $Y=52340
X14 35 M3_M2_CDNS_2 $T=78550 36430 0 0 $X=78470 $Y=36180
X15 39 M3_M2_CDNS_2 $T=79400 52420 0 90 $X=79150 $Y=52340
X16 36 M3_M2_CDNS_2 $T=86760 34460 0 0 $X=86680 $Y=34210
X17 37 M3_M2_CDNS_2 $T=86760 49100 0 0 $X=86680 $Y=48850
X18 35 M2_M1_CDNS_3 $T=51080 34160 0 0 $X=51000 $Y=33910
X19 2 M2_M1_CDNS_3 $T=52330 32180 0 90 $X=52080 $Y=32100
X20 35 M2_M1_CDNS_3 $T=52330 46820 0 90 $X=52080 $Y=46740
X21 40 M2_M1_CDNS_3 $T=54270 29810 0 90 $X=54020 $Y=29730
X22 41 M2_M1_CDNS_3 $T=54270 44450 0 90 $X=54020 $Y=44370
X23 42 M2_M1_CDNS_3 $T=55540 26280 0 0 $X=55460 $Y=26030
X24 43 M2_M1_CDNS_3 $T=55540 40920 0 0 $X=55460 $Y=40670
X25 44 M2_M1_CDNS_3 $T=55730 21200 0 90 $X=55480 $Y=21120
X26 45 M2_M1_CDNS_3 $T=55730 35840 0 90 $X=55480 $Y=35760
X27 46 M2_M1_CDNS_3 $T=56210 23810 0 90 $X=55960 $Y=23730
X28 47 M2_M1_CDNS_3 $T=56210 38450 0 90 $X=55960 $Y=38370
X29 48 M2_M1_CDNS_3 $T=56050 31070 0 0 $X=55970 $Y=30820
X30 49 M2_M1_CDNS_3 $T=56050 45710 0 0 $X=55970 $Y=45460
X31 36 M2_M1_CDNS_3 $T=56340 32800 0 0 $X=56260 $Y=32550
X32 37 M2_M1_CDNS_3 $T=56340 47440 0 0 $X=56260 $Y=47190
X33 38 M2_M1_CDNS_3 $T=57240 50840 0 0 $X=57160 $Y=50590
X34 13 M2_M1_CDNS_3 $T=57660 26200 0 90 $X=57410 $Y=26120
X35 11 M2_M1_CDNS_3 $T=57660 33520 0 90 $X=57410 $Y=33440
X36 10 M2_M1_CDNS_3 $T=57660 40840 0 90 $X=57410 $Y=40760
X37 8 M2_M1_CDNS_3 $T=57660 48160 0 90 $X=57410 $Y=48080
X38 7 M2_M1_CDNS_3 $T=57670 22770 0 90 $X=57420 $Y=22690
X39 12 M2_M1_CDNS_3 $T=57670 30070 0 90 $X=57420 $Y=29990
X40 6 M2_M1_CDNS_3 $T=57670 37410 0 90 $X=57420 $Y=37330
X41 9 M2_M1_CDNS_3 $T=57670 44710 0 90 $X=57420 $Y=44630
X42 39 M2_M1_CDNS_3 $T=72650 52420 0 90 $X=72400 $Y=52340
X43 35 M2_M1_CDNS_3 $T=78550 36430 0 0 $X=78470 $Y=36180
X44 39 M2_M1_CDNS_3 $T=79400 52420 0 90 $X=79150 $Y=52340
X45 36 M2_M1_CDNS_3 $T=86760 34460 0 0 $X=86680 $Y=34210
X46 37 M2_M1_CDNS_3 $T=86760 49100 0 0 $X=86680 $Y=48850
X47 2 M1_PO_CDNS_6 $T=52330 32180 0 90 $X=52080 $Y=32080
X48 35 M1_PO_CDNS_6 $T=52330 46820 0 90 $X=52080 $Y=46720
X49 40 M1_PO_CDNS_6 $T=54270 29810 0 90 $X=54020 $Y=29710
X50 41 M1_PO_CDNS_6 $T=54270 44450 0 90 $X=54020 $Y=44350
X51 42 M1_PO_CDNS_6 $T=55540 26280 0 0 $X=55440 $Y=26030
X52 43 M1_PO_CDNS_6 $T=55540 40920 0 0 $X=55440 $Y=40670
X53 44 M1_PO_CDNS_6 $T=55730 21200 0 90 $X=55480 $Y=21100
X54 45 M1_PO_CDNS_6 $T=55730 35840 0 90 $X=55480 $Y=35740
X55 48 M1_PO_CDNS_6 $T=56050 31070 0 0 $X=55950 $Y=30820
X56 49 M1_PO_CDNS_6 $T=56050 45710 0 0 $X=55950 $Y=45460
X57 46 M1_PO_CDNS_6 $T=56210 23810 0 90 $X=55960 $Y=23710
X58 47 M1_PO_CDNS_6 $T=56210 38450 0 90 $X=55960 $Y=38350
X59 36 M1_PO_CDNS_6 $T=56340 32800 0 0 $X=56240 $Y=32550
X60 37 M1_PO_CDNS_6 $T=56340 47440 0 0 $X=56240 $Y=47190
X61 13 M1_PO_CDNS_6 $T=57660 26200 0 90 $X=57410 $Y=26100
X62 11 M1_PO_CDNS_6 $T=57660 33520 0 90 $X=57410 $Y=33420
X63 10 M1_PO_CDNS_6 $T=57660 40840 0 90 $X=57410 $Y=40740
X64 8 M1_PO_CDNS_6 $T=57660 48160 0 90 $X=57410 $Y=48060
X65 7 M1_PO_CDNS_6 $T=57670 22770 0 90 $X=57420 $Y=22670
X66 12 M1_PO_CDNS_6 $T=57670 30070 0 90 $X=57420 $Y=29970
X67 6 M1_PO_CDNS_6 $T=57670 37410 0 90 $X=57420 $Y=37310
X68 9 M1_PO_CDNS_6 $T=57670 44710 0 90 $X=57420 $Y=44610
X69 35 M1_PO_CDNS_6 $T=78550 36430 0 0 $X=78450 $Y=36180
X70 3 M2_M1_CDNS_8 $T=50480 50560 0 0 $X=50400 $Y=50430
X71 3 M2_M1_CDNS_8 $T=51590 45750 0 90 $X=51460 $Y=45670
X72 50 M2_M1_CDNS_8 $T=53210 27000 0 0 $X=53130 $Y=26870
X73 51 M2_M1_CDNS_8 $T=53210 41640 0 0 $X=53130 $Y=41510
X74 52 M2_M1_CDNS_8 $T=53230 23140 0 0 $X=53150 $Y=23010
X75 53 M2_M1_CDNS_8 $T=53230 37780 0 0 $X=53150 $Y=37650
X76 3 M2_M1_CDNS_8 $T=62920 24380 0 0 $X=62840 $Y=24250
X77 3 M2_M1_CDNS_8 $T=62920 39020 0 0 $X=62840 $Y=38890
X78 3 M2_M1_CDNS_8 $T=62930 31710 0 0 $X=62850 $Y=31580
X79 3 M2_M1_CDNS_8 $T=62930 46350 0 0 $X=62850 $Y=46220
X80 2 M3_M2_CDNS_9 $T=52330 32180 0 90 $X=52080 $Y=32100
X81 35 M3_M2_CDNS_9 $T=52330 46820 0 90 $X=52080 $Y=46740
X82 42 M3_M2_CDNS_9 $T=53480 29020 0 0 $X=53400 $Y=28770
X83 43 M3_M2_CDNS_9 $T=53480 43660 0 0 $X=53400 $Y=43410
X84 40 M3_M2_CDNS_9 $T=54270 29810 0 90 $X=54020 $Y=29730
X85 41 M3_M2_CDNS_9 $T=54270 44450 0 90 $X=54020 $Y=44370
X86 42 M3_M2_CDNS_9 $T=55540 26280 0 0 $X=55460 $Y=26030
X87 43 M3_M2_CDNS_9 $T=55540 40920 0 0 $X=55460 $Y=40670
X88 44 M3_M2_CDNS_9 $T=55730 21200 0 90 $X=55480 $Y=21120
X89 45 M3_M2_CDNS_9 $T=55730 35840 0 90 $X=55480 $Y=35760
X90 46 M3_M2_CDNS_9 $T=56210 23810 0 90 $X=55960 $Y=23730
X91 47 M3_M2_CDNS_9 $T=56210 38450 0 90 $X=55960 $Y=38370
X92 48 M3_M2_CDNS_9 $T=56050 31070 0 0 $X=55970 $Y=30820
X93 49 M3_M2_CDNS_9 $T=56050 45710 0 0 $X=55970 $Y=45460
X94 50 M3_M2_CDNS_9 $T=56240 34220 0 0 $X=56160 $Y=33970
X95 51 M3_M2_CDNS_9 $T=56240 48860 0 0 $X=56160 $Y=48610
X96 13 M3_M2_CDNS_9 $T=57660 26200 0 90 $X=57410 $Y=26120
X97 11 M3_M2_CDNS_9 $T=57660 33520 0 90 $X=57410 $Y=33440
X98 10 M3_M2_CDNS_9 $T=57660 40840 0 90 $X=57410 $Y=40760
X99 8 M3_M2_CDNS_9 $T=57660 48160 0 90 $X=57410 $Y=48080
X100 7 M3_M2_CDNS_9 $T=57670 22770 0 90 $X=57420 $Y=22690
X101 12 M3_M2_CDNS_9 $T=57670 30070 0 90 $X=57420 $Y=29990
X102 6 M3_M2_CDNS_9 $T=57670 37410 0 90 $X=57420 $Y=37330
X103 9 M3_M2_CDNS_9 $T=57670 44710 0 90 $X=57420 $Y=44630
X104 48 M3_M2_CDNS_9 $T=62950 31240 0 90 $X=62700 $Y=31160
X105 49 M3_M2_CDNS_9 $T=62950 45880 0 90 $X=62700 $Y=45800
X106 46 M3_M2_CDNS_9 $T=63400 23460 0 0 $X=63320 $Y=23210
X107 47 M3_M2_CDNS_9 $T=63400 38100 0 0 $X=63320 $Y=37850
X108 44 M3_M2_CDNS_9 $T=63720 21760 0 0 $X=63640 $Y=21510
X109 45 M3_M2_CDNS_9 $T=63720 36400 0 0 $X=63640 $Y=36150
X110 40 M3_M2_CDNS_9 $T=63820 29420 0 0 $X=63740 $Y=29170
X111 41 M3_M2_CDNS_9 $T=63820 44060 0 0 $X=63740 $Y=43810
X112 50 M3_M2_CDNS_10 $T=50730 34460 0 0 $X=50650 $Y=34330
X113 51 M3_M2_CDNS_10 $T=50800 49100 0 0 $X=50720 $Y=48970
X114 2 M3_M2_CDNS_10 $T=51610 22610 0 0 $X=51530 $Y=22480
X115 35 M4_M3_CDNS_12 $T=51140 36930 0 0 $X=51060 $Y=36800
X116 42 M2_M1_CDNS_13 $T=53480 29020 0 0 $X=53400 $Y=28770
X117 43 M2_M1_CDNS_13 $T=53480 43660 0 0 $X=53400 $Y=43410
X118 50 M2_M1_CDNS_13 $T=56240 34220 0 0 $X=56160 $Y=33970
X119 51 M2_M1_CDNS_13 $T=56240 48860 0 0 $X=56160 $Y=48610
X120 48 M2_M1_CDNS_13 $T=62950 31240 0 90 $X=62700 $Y=31160
X121 49 M2_M1_CDNS_13 $T=62950 45880 0 90 $X=62700 $Y=45800
X122 46 M2_M1_CDNS_13 $T=63400 23460 0 0 $X=63320 $Y=23210
X123 47 M2_M1_CDNS_13 $T=63400 38100 0 0 $X=63320 $Y=37850
X124 44 M2_M1_CDNS_13 $T=63720 21760 0 0 $X=63640 $Y=21510
X125 45 M2_M1_CDNS_13 $T=63720 36400 0 0 $X=63640 $Y=36150
X126 40 M2_M1_CDNS_13 $T=63820 29420 0 0 $X=63740 $Y=29170
X127 41 M2_M1_CDNS_13 $T=63820 44060 0 0 $X=63740 $Y=43810
X128 52 M1_PO_CDNS_15 $T=53520 24980 0 90 $X=53270 $Y=24880
X129 53 M1_PO_CDNS_15 $T=53520 39620 0 90 $X=53270 $Y=39520
X130 14 M1_PO_CDNS_15 $T=64110 23330 0 0 $X=64010 $Y=23080
X131 18 M1_PO_CDNS_15 $T=64110 37970 0 0 $X=64010 $Y=37720
X132 14 M1_PO_CDNS_15 $T=65950 23850 0 90 $X=65700 $Y=23750
X133 18 M1_PO_CDNS_15 $T=65950 38490 0 90 $X=65700 $Y=38390
X134 2 M1_PO_CDNS_15 $T=78510 22370 0 0 $X=78410 $Y=22120
X135 54 M1_PO_CDNS_16 $T=53270 31100 0 0 $X=53170 $Y=30980
X136 55 M1_PO_CDNS_16 $T=53270 45740 0 0 $X=53170 $Y=45620
X137 56 M1_PO_CDNS_16 $T=53550 23450 0 0 $X=53450 $Y=23330
X138 57 M1_PO_CDNS_16 $T=53550 38090 0 0 $X=53450 $Y=37970
X139 58 M1_PO_CDNS_16 $T=53840 25910 0 0 $X=53740 $Y=25790
X140 59 M1_PO_CDNS_16 $T=53840 40550 0 0 $X=53740 $Y=40430
X141 52 M2_M1_CDNS_17 $T=53520 24980 0 90 $X=53270 $Y=24900
X142 53 M2_M1_CDNS_17 $T=53520 39620 0 90 $X=53270 $Y=39540
X143 14 M2_M1_CDNS_17 $T=64110 23330 0 0 $X=64030 $Y=23080
X144 18 M2_M1_CDNS_17 $T=64110 37970 0 0 $X=64030 $Y=37720
X145 14 M2_M1_CDNS_17 $T=65950 23850 0 90 $X=65700 $Y=23770
X146 18 M2_M1_CDNS_17 $T=65950 38490 0 90 $X=65700 $Y=38410
X147 2 M2_M1_CDNS_17 $T=78510 22370 0 0 $X=78430 $Y=22120
X148 3 4 44 56 46 172 NAND_1X_small $T=53960 20720 0 0 $X=53530 $Y=20700
X149 3 4 42 58 52 171 NAND_1X_small $T=55940 28040 0 180 $X=53530 $Y=24260
X150 3 4 40 54 48 170 NAND_1X_small $T=53960 28040 0 0 $X=53530 $Y=28020
X151 3 4 45 57 47 169 NAND_1X_small $T=53960 35360 0 0 $X=53530 $Y=35340
X152 3 4 43 59 53 168 NAND_1X_small $T=55940 42680 0 180 $X=53530 $Y=38900
X153 3 4 41 55 49 167 NAND_1X_small $T=53960 42680 0 0 $X=53530 $Y=42660
X154 3 4 14 7 46 85 86 187 265 188 XOR1 $T=56070 20720 0 0 $X=56130 $Y=20700
X155 3 4 15 13 44 83 84 185 264 186 XOR1 $T=56070 28040 1 0 $X=56130 $Y=24260
X156 3 4 16 12 48 81 82 183 263 184 XOR1 $T=56070 28040 0 0 $X=56130 $Y=28020
X157 3 4 17 11 40 79 80 181 262 182 XOR1 $T=56070 35360 1 0 $X=56130 $Y=31580
X158 3 4 18 6 47 77 78 179 261 180 XOR1 $T=56070 35360 0 0 $X=56130 $Y=35340
X159 3 4 19 10 45 75 76 177 260 178 XOR1 $T=56070 42680 1 0 $X=56130 $Y=38900
X160 3 4 20 9 49 73 74 175 259 176 XOR1 $T=56070 42680 0 0 $X=56130 $Y=42660
X161 3 4 21 8 41 71 72 173 258 174 XOR1 $T=56070 50000 1 0 $X=56130 $Y=46220
X162 5 3 1 4 38 22 39 66 69 70
+ 64 65 67 68 256 257 full_adder1_small $T=50650 49970 0 0 $X=50670 $Y=49980
X163 24 3 23 4 39 33 34 151 154 155
+ 149 150 152 153 266 267 full_adder1_small $T=72610 49970 0 0 $X=72630 $Y=49980
X164 50 36 3 4 2 35 62 63 158 159
+ 254 255 MUX_2to1___2X $T=56190 30160 0 180 $X=50640 $Y=31580
X165 51 37 3 4 35 38 60 61 156 157
+ 252 253 MUX_2to1___2X $T=56190 44800 0 180 $X=50640 $Y=46220
X166 14 13 12 11 3 7 4 15 16 17
+ 2 25 28 27 26 36 138 139 140 FA_4bit $T=64900 20820 0 0 $X=64250 $Y=20700
X167 18 10 9 8 3 6 4 19 20 21
+ 35 32 31 30 29 37 107 108 109 FA_4bit $T=64900 35460 0 0 $X=64250 $Y=35340
X168 56 3 4 52 INV_1X_small $T=51530 20700 0 0 $X=51530 $Y=20700
X169 58 3 4 50 INV_1X_small $T=51530 28060 1 0 $X=51530 $Y=24260
X170 54 3 4 42 INV_1X_small $T=51530 28020 0 0 $X=51530 $Y=28020
X171 57 3 4 53 INV_1X_small $T=51530 35340 0 0 $X=51530 $Y=35340
X172 59 3 4 51 INV_1X_small $T=51530 42700 1 0 $X=51530 $Y=38900
X173 55 3 4 43 INV_1X_small $T=51530 42660 0 0 $X=51530 $Y=42660
M0 64 5 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6612 scb=0.0167915 scc=0.000377457 $X=51440 $Y=52320 $dt=1
M1 65 1 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.8911 scb=0.00996238 scc=0.000256798 $X=52400 $Y=52320 $dt=1
M2 256 1 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=53730 $Y=52080 $dt=1
M3 58 52 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=25230 $dt=1
M4 59 53 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=39870 $dt=1
M5 66 64 256 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=54700 $Y=52140 $dt=1
M6 56 44 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=23050 $dt=1
M7 54 40 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=30370 $dt=1
M8 57 45 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=37690 $dt=1
M9 55 41 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=45010 $dt=1
M10 3 42 58 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=25230 $dt=1
M11 3 43 59 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=39870 $dt=1
M12 3 46 56 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=23050 $dt=1
M13 3 48 54 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=30370 $dt=1
M14 3 47 57 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=37690 $dt=1
M15 3 49 55 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=45010 $dt=1
M16 66 65 256 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=55660 $Y=52140 $dt=1
M17 256 5 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=56620 $Y=52140 $dt=1
M18 85 14 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=23040 $dt=1
M19 83 15 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=25240 $dt=1
M20 81 16 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=30360 $dt=1
M21 79 17 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=32560 $dt=1
M22 77 18 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=37680 $dt=1
M23 75 19 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=39880 $dt=1
M24 73 20 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=45000 $dt=1
M25 71 21 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=47200 $dt=1
M26 86 7 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=23040 $dt=1
M27 84 13 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=25240 $dt=1
M28 82 12 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=30360 $dt=1
M29 80 11 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=32560 $dt=1
M30 78 6 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=37680 $dt=1
M31 76 10 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=39880 $dt=1
M32 74 9 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=45000 $dt=1
M33 72 8 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=47200 $dt=1
M34 67 38 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=58280 $Y=52320 $dt=1
M35 265 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=22800 $dt=1
M36 264 13 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=25000 $dt=1
M37 263 12 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=30120 $dt=1
M38 262 11 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=32320 $dt=1
M39 261 6 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=37440 $dt=1
M40 260 10 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=39640 $dt=1
M41 259 9 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=44760 $dt=1
M42 258 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=46960 $dt=1
M43 68 66 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=59240 $Y=52320 $dt=1
M44 46 85 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=22860 $dt=1
M45 44 83 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=24940 $dt=1
M46 48 81 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=30180 $dt=1
M47 40 79 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=32260 $dt=1
M48 47 77 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=37500 $dt=1
M49 45 75 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=39580 $dt=1
M50 49 73 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=44820 $dt=1
M51 41 71 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=46900 $dt=1
M52 257 66 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60570 $Y=52080 $dt=1
M53 46 86 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=22860 $dt=1
M54 44 84 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=24940 $dt=1
M55 48 82 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=30180 $dt=1
M56 40 80 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=32260 $dt=1
M57 47 78 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=37500 $dt=1
M58 45 76 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=39580 $dt=1
M59 49 74 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=44820 $dt=1
M60 41 72 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=46900 $dt=1
M61 22 67 257 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=61540 $Y=52140 $dt=1
M62 265 14 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=22860 $dt=1
M63 264 15 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=24940 $dt=1
M64 263 16 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=30180 $dt=1
M65 262 17 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=32260 $dt=1
M66 261 18 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=37500 $dt=1
M67 260 19 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=39580 $dt=1
M68 259 20 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=44820 $dt=1
M69 258 21 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=46900 $dt=1
M70 22 68 257 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=62500 $Y=52140 $dt=1
M71 257 38 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=63460 $Y=52140 $dt=1
M72 69 38 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65530 $Y=52110 $dt=1
M73 3 66 69 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65940 $Y=52110 $dt=1
M74 70 5 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68510 $Y=52330 $dt=1
M75 3 1 70 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68920 $Y=52330 $dt=1
M76 39 69 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71350 $Y=52330 $dt=1
M77 3 70 39 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71760 $Y=52330 $dt=1
M78 149 24 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=73400 $Y=52320 $dt=1
M79 150 23 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=74360 $Y=52320 $dt=1
M80 266 23 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=75690 $Y=52080 $dt=1
M81 151 149 266 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=76660 $Y=52140 $dt=1
M82 151 150 266 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=77620 $Y=52140 $dt=1
M83 266 24 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=78580 $Y=52140 $dt=1
M84 152 39 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=80240 $Y=52320 $dt=1
M85 153 151 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=81200 $Y=52320 $dt=1
M86 267 151 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=82530 $Y=52080 $dt=1
M87 33 152 267 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=83500 $Y=52140 $dt=1
M88 33 153 267 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=84460 $Y=52140 $dt=1
M89 267 39 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=85420 $Y=52140 $dt=1
M90 154 39 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87490 $Y=52110 $dt=1
M91 3 151 154 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87900 $Y=52110 $dt=1
M92 155 24 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90470 $Y=52330 $dt=1
M93 3 23 155 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90880 $Y=52330 $dt=1
M94 34 154 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=93310 $Y=52330 $dt=1
M95 3 155 34 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=93720 $Y=52330 $dt=1
.ends 10badder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_46                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_46 1 2 3 5
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=660 $Y=760 $dt=0
.ends cellTmpl_CDNS_46

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 1 M1_PO_CDNS_16 $T=700 2040 0 90 $X=580 $Y=1940
X1 2 3 1 4 cellTmpl_CDNS_46 $T=120 140 0 0 $X=0 $Y=0
.ends INV_1X_small_layout

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_16 $T=640 1830 0 90 $X=520 $Y=1730
X1 6 M1_PO_CDNS_16 $T=1940 640 0 0 $X=1840 $Y=520
X2 3 1 6 3 nmos1v_CDNS_19 $T=710 860 0 0 $X=290 $Y=660
X3 4 6 5 3 nmos1v_CDNS_19 $T=1890 860 0 0 $X=1470 $Y=660
X4 2 3 cellTmpl_CDNS_21 $T=120 140 0 0 $X=0 $Y=0
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=710 $Y=860 $dt=0
M1 5 6 4 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1890 $Y=860 $dt=0
.ends ph1p3_clk_part

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_48                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_48 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_48

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_MSDFF                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_MSDFF 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17
*.DEVICECLIMB
** N=18 EP=17 FDC=15
X0 1 M4_M3_CDNS_1 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X1 1 M4_M3_CDNS_1 $T=5110 3310 0 0 $X=5030 $Y=3060
X2 1 M3_M2_CDNS_2 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X3 1 M3_M2_CDNS_2 $T=5110 3310 0 0 $X=5030 $Y=3060
X4 1 M2_M1_CDNS_3 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X5 1 M2_M1_CDNS_3 $T=5110 3310 0 0 $X=5030 $Y=3060
X6 7 M2_M1_CDNS_3 $T=8100 2170 0 90 $X=7850 $Y=2090
X7 7 M1_PO_CDNS_6 $T=8100 2170 0 90 $X=7850 $Y=2070
X8 2 M2_M1_CDNS_8 $T=430 2010 0 0 $X=350 $Y=1880
X9 8 M2_M1_CDNS_8 $T=1110 -1470 0 0 $X=1030 $Y=-1600
X10 2 M2_M1_CDNS_8 $T=2790 -1820 0 0 $X=2710 $Y=-1950
X11 9 M2_M1_CDNS_8 $T=4150 -1460 0 0 $X=4070 $Y=-1590
X12 6 M2_M1_CDNS_8 $T=5200 -2030 0 0 $X=5120 $Y=-2160
X13 8 M2_M1_CDNS_8 $T=5310 1560 0 90 $X=5180 $Y=1480
X14 9 M2_M1_CDNS_8 $T=5670 -1460 0 90 $X=5540 $Y=-1540
X15 10 M2_M1_CDNS_8 $T=6280 1490 0 0 $X=6200 $Y=1360
X16 11 M2_M1_CDNS_8 $T=7300 1510 0 90 $X=7170 $Y=1430
X17 10 M2_M1_CDNS_8 $T=7850 -2080 0 0 $X=7770 $Y=-2210
X18 11 M2_M1_CDNS_8 $T=9400 1510 0 90 $X=9270 $Y=1430
X19 6 M2_M1_CDNS_8 $T=9770 -2060 0 0 $X=9690 $Y=-2190
X20 7 M3_M2_CDNS_9 $T=1140 2170 0 90 $X=890 $Y=2090
X21 12 M3_M2_CDNS_9 $T=3910 970 0 0 $X=3830 $Y=720
X22 13 M3_M2_CDNS_9 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X23 7 M3_M2_CDNS_9 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X24 7 M3_M2_CDNS_9 $T=8100 2170 0 90 $X=7850 $Y=2090
X25 13 M3_M2_CDNS_9 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X26 12 M3_M2_CDNS_9 $T=9760 1890 0 0 $X=9680 $Y=1640
X27 7 M2_M1_CDNS_13 $T=1140 2170 0 90 $X=890 $Y=2090
X28 12 M2_M1_CDNS_13 $T=3910 970 0 0 $X=3830 $Y=720
X29 13 M2_M1_CDNS_13 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X30 7 M2_M1_CDNS_13 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X31 13 M2_M1_CDNS_13 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X32 12 M2_M1_CDNS_13 $T=9760 1890 0 0 $X=9680 $Y=1640
X33 12 1 3 8 10 18 NAND2_1X_small $T=3680 -70 0 0 $X=3800 $Y=0
X34 4 1 3 8 INV_1X_small_layout $T=0 40 1 0 $X=0 $Y=-3760
X35 2 1 3 7 INV_1X_small_layout $T=0 0 0 0 $X=0 $Y=0
X36 6 1 3 9 INV_1X_small_layout $T=4800 40 1 0 $X=4800 $Y=-3760
X37 10 1 3 11 INV_1X_small_layout $T=6200 0 0 0 $X=6200 $Y=0
X38 13 1 3 6 INV_1X_small_layout $T=8600 40 1 0 $X=8600 $Y=-3760
X39 2 1 3 5 12 14 ph1p3_clk_part $T=1400 0 0 0 $X=1400 $Y=0
X40 2 1 3 9 13 15 ph1p3_clk_part $T=2400 40 1 0 $X=2400 $Y=-3760
X41 7 1 3 10 13 16 ph1p3_clk_part $T=6200 40 1 0 $X=6200 $Y=-3760
X42 7 1 3 11 12 17 ph1p3_clk_part $T=7600 0 0 0 $X=7600 $Y=0
X43 1 3 cellTmpl_CDNS_48 $T=1520 -100 1 0 $X=1400 $Y=-3760
.ends ph1p3_MSDFF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_49                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_49 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_49

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X_ph2p2                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X_ph2p2 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=12 EP=12 FDC=6
X0 7 M2_M1_CDNS_3 $T=430 2220 0 0 $X=350 $Y=1970
X1 7 M2_M1_CDNS_3 $T=2800 2490 0 0 $X=2720 $Y=2240
X2 7 M1_PO_CDNS_6 $T=430 2220 0 0 $X=330 $Y=1970
X3 7 M1_PO_CDNS_6 $T=2800 2490 0 0 $X=2700 $Y=2240
X4 7 M3_M2_CDNS_9 $T=430 2220 0 0 $X=350 $Y=1970
X5 7 M3_M2_CDNS_9 $T=1140 3180 0 0 $X=1060 $Y=2930
X6 7 M3_M2_CDNS_9 $T=2800 2490 0 0 $X=2720 $Y=2240
X7 7 M2_M1_CDNS_13 $T=1140 3180 0 0 $X=1060 $Y=2930
X8 1 M1_PO_CDNS_15 $T=1480 1720 0 0 $X=1380 $Y=1470
X9 1 M1_PO_CDNS_15 $T=2840 980 0 0 $X=2740 $Y=730
X10 1 M1_PO_CDNS_16 $T=860 1670 0 0 $X=760 $Y=1550
X11 2 M1_PO_CDNS_16 $T=1480 3130 0 0 $X=1380 $Y=3010
X12 5 M1_PO_CDNS_16 $T=4220 2040 0 0 $X=4120 $Y=1920
X13 8 M1_PO_CDNS_16 $T=4480 1550 0 90 $X=4360 $Y=1450
X14 1 M2_M1_CDNS_17 $T=1480 1720 0 0 $X=1400 $Y=1470
X15 1 M2_M1_CDNS_17 $T=2840 980 0 0 $X=2760 $Y=730
X16 4 7 9 4 nmos1v_CDNS_31 $T=2170 800 0 0 $X=1970 $Y=600
X17 8 5 10 4 nmos1v_CDNS_31 $T=3550 790 0 0 $X=3350 $Y=590
X18 8 2 9 4 nmos1v_CDNS_32 $T=1960 800 0 0 $X=1540 $Y=600
X19 4 1 10 4 nmos1v_CDNS_32 $T=3340 790 0 0 $X=2920 $Y=590
X20 3 4 1 7 8 6 cellTmpl_CDNS_43 $T=120 140 0 0 $X=0 $Y=0
X21 3 1 11 4 3 pmos1v_CDNS_44 $T=2170 2100 0 0 $X=1970 $Y=1900
X22 8 5 12 4 3 pmos1v_CDNS_44 $T=3550 2030 0 0 $X=3350 $Y=1830
X23 8 2 11 4 3 pmos1v_CDNS_45 $T=1960 2100 0 0 $X=1540 $Y=1900
X24 3 7 12 4 3 pmos1v_CDNS_45 $T=3340 2030 0 0 $X=2920 $Y=1830
M0 9 2 8 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1960 $Y=800 $dt=0
M1 4 7 9 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=2170 $Y=800 $dt=0
M2 10 1 4 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3340 $Y=790 $dt=0
M3 8 5 10 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3550 $Y=790 $dt=0
.ends MUX_2to1___2X_ph2p2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p2_processing_element                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p2_processing_element 26 24 23 18 43 44 52 50 48 46
+ 21 22 20 19 47 49 51 53 15 42
+ 33 54 17 73 71 69 67 63 59 55
+ 65 61 57 74 72 70 68 64 60 56
+ 66 62 58 1 41
** N=785 EP=45 FDC=1662
X0 1 M4_M3_CDNS_1 $T=1340 55390 0 0 $X=1260 $Y=55140
X1 1 M4_M3_CDNS_1 $T=3450 61970 0 0 $X=3370 $Y=61720
X2 1 M4_M3_CDNS_1 $T=9870 69280 0 0 $X=9790 $Y=69030
X3 2 M4_M3_CDNS_1 $T=14700 34240 0 0 $X=14620 $Y=33990
X4 3 M4_M3_CDNS_1 $T=15150 34320 0 0 $X=15070 $Y=34070
X5 4 M4_M3_CDNS_1 $T=28040 20980 0 0 $X=27960 $Y=20730
X6 5 M4_M3_CDNS_1 $T=30360 48950 0 0 $X=30280 $Y=48700
X7 6 M4_M3_CDNS_1 $T=30540 30290 0 90 $X=30290 $Y=30210
X8 7 M4_M3_CDNS_1 $T=30920 28440 0 90 $X=30670 $Y=28360
X9 7 M4_M3_CDNS_1 $T=30920 23090 0 0 $X=30840 $Y=22840
X10 6 M4_M3_CDNS_1 $T=30960 32190 0 0 $X=30880 $Y=31940
X11 8 M4_M3_CDNS_1 $T=34240 15510 0 0 $X=34160 $Y=15260
X12 9 M4_M3_CDNS_1 $T=36070 26280 0 0 $X=35990 $Y=26030
X13 6 M4_M3_CDNS_1 $T=36600 41550 0 0 $X=36520 $Y=41300
X14 10 M4_M3_CDNS_1 $T=37620 30320 0 0 $X=37540 $Y=30070
X15 11 M4_M3_CDNS_1 $T=37800 29000 0 0 $X=37720 $Y=28750
X16 6 M4_M3_CDNS_1 $T=38820 45300 0 0 $X=38740 $Y=45050
X17 12 M4_M3_CDNS_1 $T=40600 12040 0 0 $X=40520 $Y=11790
X18 12 M4_M3_CDNS_1 $T=40600 13810 0 0 $X=40520 $Y=13560
X19 13 M4_M3_CDNS_1 $T=41660 8130 0 0 $X=41580 $Y=7880
X20 14 M4_M3_CDNS_1 $T=43120 8620 0 0 $X=43040 $Y=8370
X21 15 M4_M3_CDNS_1 $T=45720 13840 0 0 $X=45640 $Y=13590
X22 15 M4_M3_CDNS_1 $T=46890 13630 0 0 $X=46810 $Y=13380
X23 15 M4_M3_CDNS_1 $T=46900 20740 0 0 $X=46820 $Y=20490
X24 15 M4_M3_CDNS_1 $T=46910 28080 0 0 $X=46830 $Y=27830
X25 1 M4_M3_CDNS_1 $T=49180 4060 0 0 $X=49100 $Y=3810
X26 1 M4_M3_CDNS_1 $T=49180 11470 0 0 $X=49100 $Y=11220
X27 1 M4_M3_CDNS_1 $T=49180 18800 0 0 $X=49100 $Y=18550
X28 1 M4_M3_CDNS_1 $T=49180 26120 0 0 $X=49100 $Y=25870
X29 1 M4_M3_CDNS_1 $T=49180 33430 0 0 $X=49100 $Y=33180
X30 1 M4_M3_CDNS_1 $T=49180 40820 0 0 $X=49100 $Y=40570
X31 1 M4_M3_CDNS_1 $T=49180 48070 0 0 $X=49100 $Y=47820
X32 1 M4_M3_CDNS_1 $T=49180 54710 0 0 $X=49100 $Y=54460
X33 16 M4_M3_CDNS_1 $T=50830 40760 0 90 $X=50580 $Y=40680
X34 17 M4_M3_CDNS_1 $T=58260 1650 0 0 $X=58180 $Y=1400
X35 17 M4_M3_CDNS_1 $T=58670 9650 0 90 $X=58420 $Y=9570
X36 17 M4_M3_CDNS_1 $T=58670 12550 0 90 $X=58420 $Y=12470
X37 17 M4_M3_CDNS_1 $T=58670 16970 0 90 $X=58420 $Y=16890
X38 17 M4_M3_CDNS_1 $T=58670 19870 0 90 $X=58420 $Y=19790
X39 17 M4_M3_CDNS_1 $T=58670 24290 0 90 $X=58420 $Y=24210
X40 17 M4_M3_CDNS_1 $T=58670 27190 0 90 $X=58420 $Y=27110
X41 17 M4_M3_CDNS_1 $T=58670 31610 0 90 $X=58420 $Y=31530
X42 17 M4_M3_CDNS_1 $T=58670 38930 0 90 $X=58420 $Y=38850
X43 17 M4_M3_CDNS_1 $T=58670 46250 0 90 $X=58420 $Y=46170
X44 17 M4_M3_CDNS_1 $T=58670 53570 0 90 $X=58420 $Y=53490
X45 1 M3_M2_CDNS_2 $T=1340 55390 0 0 $X=1260 $Y=55140
X46 18 M3_M2_CDNS_2 $T=1480 56760 0 0 $X=1400 $Y=56510
X47 19 M3_M2_CDNS_2 $T=2350 44590 0 90 $X=2100 $Y=44510
X48 1 M3_M2_CDNS_2 $T=3450 61970 0 0 $X=3370 $Y=61720
X49 20 M3_M2_CDNS_2 $T=3900 48300 0 90 $X=3650 $Y=48220
X50 21 M3_M2_CDNS_2 $T=3940 58210 0 90 $X=3690 $Y=58130
X51 18 M3_M2_CDNS_2 $T=4250 65060 0 180 $X=4170 $Y=64810
X52 21 M3_M2_CDNS_2 $T=4250 72470 0 0 $X=4170 $Y=72220
X53 22 M3_M2_CDNS_2 $T=6840 58120 0 90 $X=6590 $Y=58040
X54 1 M3_M2_CDNS_2 $T=9870 69280 0 0 $X=9790 $Y=69030
X55 23 M3_M2_CDNS_2 $T=11380 56560 0 90 $X=11130 $Y=56480
X56 23 M3_M2_CDNS_2 $T=14490 65150 0 0 $X=14410 $Y=64900
X57 22 M3_M2_CDNS_2 $T=14490 72480 0 0 $X=14410 $Y=72230
X58 2 M3_M2_CDNS_2 $T=14700 34240 0 0 $X=14620 $Y=33990
X59 24 M3_M2_CDNS_2 $T=20420 56560 0 90 $X=20170 $Y=56480
X60 24 M3_M2_CDNS_2 $T=24730 65150 0 0 $X=24650 $Y=64900
X61 20 M3_M2_CDNS_2 $T=24730 72470 0 0 $X=24650 $Y=72220
X62 25 M3_M2_CDNS_2 $T=27620 26990 0 0 $X=27540 $Y=26740
X63 4 M3_M2_CDNS_2 $T=28040 20980 0 0 $X=27960 $Y=20730
X64 26 M3_M2_CDNS_2 $T=29230 56560 0 90 $X=28980 $Y=56480
X65 27 M3_M2_CDNS_2 $T=32470 34080 0 90 $X=32220 $Y=34000
X66 28 M3_M2_CDNS_2 $T=33670 6150 0 90 $X=33420 $Y=6070
X67 26 M3_M2_CDNS_2 $T=34970 65150 0 0 $X=34890 $Y=64900
X68 19 M3_M2_CDNS_2 $T=34970 72470 0 0 $X=34890 $Y=72220
X69 29 M3_M2_CDNS_2 $T=35130 53970 0 0 $X=35050 $Y=53720
X70 10 M3_M2_CDNS_2 $T=37620 30320 0 0 $X=37540 $Y=30070
X71 30 M3_M2_CDNS_2 $T=38220 15840 0 0 $X=38140 $Y=15590
X72 28 M3_M2_CDNS_2 $T=38250 22590 0 0 $X=38170 $Y=22340
X73 31 M3_M2_CDNS_2 $T=38270 21170 0 0 $X=38190 $Y=20920
X74 6 M3_M2_CDNS_2 $T=38820 45300 0 0 $X=38740 $Y=45050
X75 12 M3_M2_CDNS_2 $T=40600 13810 0 0 $X=40520 $Y=13560
X76 32 M3_M2_CDNS_2 $T=40710 21060 0 0 $X=40630 $Y=20810
X77 15 M3_M2_CDNS_2 $T=46890 13630 0 0 $X=46810 $Y=13380
X78 15 M3_M2_CDNS_2 $T=46900 20740 0 0 $X=46820 $Y=20490
X79 15 M3_M2_CDNS_2 $T=46910 28080 0 0 $X=46830 $Y=27830
X80 14 M3_M2_CDNS_2 $T=47280 7640 0 90 $X=47030 $Y=7560
X81 30 M3_M2_CDNS_2 $T=47850 15290 0 0 $X=47770 $Y=15040
X82 28 M3_M2_CDNS_2 $T=47850 23870 0 0 $X=47770 $Y=23620
X83 33 M3_M2_CDNS_2 $T=47980 9490 0 180 $X=47900 $Y=9240
X84 33 M3_M2_CDNS_2 $T=48880 2280 0 0 $X=48800 $Y=2030
X85 1 M3_M2_CDNS_2 $T=49180 4060 0 0 $X=49100 $Y=3810
X86 1 M3_M2_CDNS_2 $T=49180 11470 0 0 $X=49100 $Y=11220
X87 1 M3_M2_CDNS_2 $T=49180 18800 0 0 $X=49100 $Y=18550
X88 1 M3_M2_CDNS_2 $T=49180 26120 0 0 $X=49100 $Y=25870
X89 1 M3_M2_CDNS_2 $T=49180 33430 0 0 $X=49100 $Y=33180
X90 1 M3_M2_CDNS_2 $T=49180 40820 0 0 $X=49100 $Y=40570
X91 1 M3_M2_CDNS_2 $T=49180 48070 0 0 $X=49100 $Y=47820
X92 1 M3_M2_CDNS_2 $T=49180 54710 0 0 $X=49100 $Y=54460
X93 15 M3_M2_CDNS_2 $T=50250 45640 0 90 $X=50000 $Y=45560
X94 13 M3_M2_CDNS_2 $T=50910 13780 0 0 $X=50830 $Y=13530
X95 17 M3_M2_CDNS_2 $T=58670 9650 0 90 $X=58420 $Y=9570
X96 17 M3_M2_CDNS_2 $T=58670 12550 0 90 $X=58420 $Y=12470
X97 17 M3_M2_CDNS_2 $T=58670 16970 0 90 $X=58420 $Y=16890
X98 17 M3_M2_CDNS_2 $T=58670 19870 0 90 $X=58420 $Y=19790
X99 17 M3_M2_CDNS_2 $T=58670 24290 0 90 $X=58420 $Y=24210
X100 17 M3_M2_CDNS_2 $T=58670 27190 0 90 $X=58420 $Y=27110
X101 17 M3_M2_CDNS_2 $T=58670 31610 0 90 $X=58420 $Y=31530
X102 17 M3_M2_CDNS_2 $T=58670 38930 0 90 $X=58420 $Y=38850
X103 17 M3_M2_CDNS_2 $T=58670 46250 0 90 $X=58420 $Y=46170
X104 17 M3_M2_CDNS_2 $T=58670 53570 0 90 $X=58420 $Y=53490
X105 14 M3_M2_CDNS_2 $T=59660 13790 0 0 $X=59580 $Y=13540
X106 30 M3_M2_CDNS_2 $T=59660 21120 0 0 $X=59580 $Y=20870
X107 28 M3_M2_CDNS_2 $T=59660 28470 0 0 $X=59580 $Y=28220
X108 1 M2_M1_CDNS_3 $T=1340 55390 0 0 $X=1260 $Y=55140
X109 18 M2_M1_CDNS_3 $T=1480 56760 0 0 $X=1400 $Y=56510
X110 33 M2_M1_CDNS_3 $T=1860 60810 0 0 $X=1780 $Y=60560
X111 33 M2_M1_CDNS_3 $T=1870 68120 0 0 $X=1790 $Y=67870
X112 19 M2_M1_CDNS_3 $T=2350 44590 0 90 $X=2100 $Y=44510
X113 1 M2_M1_CDNS_3 $T=3450 61970 0 0 $X=3370 $Y=61720
X114 20 M2_M1_CDNS_3 $T=3900 48300 0 90 $X=3650 $Y=48220
X115 21 M2_M1_CDNS_3 $T=3940 58210 0 90 $X=3690 $Y=58130
X116 18 M2_M1_CDNS_3 $T=4250 65060 0 180 $X=4170 $Y=64810
X117 21 M2_M1_CDNS_3 $T=4250 72470 0 0 $X=4170 $Y=72220
X118 22 M2_M1_CDNS_3 $T=6840 58120 0 90 $X=6590 $Y=58040
X119 1 M2_M1_CDNS_3 $T=9870 69280 0 0 $X=9790 $Y=69030
X120 23 M2_M1_CDNS_3 $T=11380 56560 0 90 $X=11130 $Y=56480
X121 33 M2_M1_CDNS_3 $T=12100 60800 0 0 $X=12020 $Y=60550
X122 33 M2_M1_CDNS_3 $T=12100 68120 0 0 $X=12020 $Y=67870
X123 23 M2_M1_CDNS_3 $T=14490 65150 0 0 $X=14410 $Y=64900
X124 22 M2_M1_CDNS_3 $T=14490 72480 0 0 $X=14410 $Y=72230
X125 24 M2_M1_CDNS_3 $T=20420 56560 0 90 $X=20170 $Y=56480
X126 33 M2_M1_CDNS_3 $T=22340 68120 0 0 $X=22260 $Y=67870
X127 33 M2_M1_CDNS_3 $T=22350 60800 0 0 $X=22270 $Y=60550
X128 24 M2_M1_CDNS_3 $T=24730 65150 0 0 $X=24650 $Y=64900
X129 20 M2_M1_CDNS_3 $T=24730 72470 0 0 $X=24650 $Y=72220
X130 25 M2_M1_CDNS_3 $T=27620 26990 0 0 $X=27540 $Y=26740
X131 4 M2_M1_CDNS_3 $T=28040 20980 0 0 $X=27960 $Y=20730
X132 26 M2_M1_CDNS_3 $T=29230 56560 0 90 $X=28980 $Y=56480
X133 33 M2_M1_CDNS_3 $T=32580 60800 0 0 $X=32500 $Y=60550
X134 33 M2_M1_CDNS_3 $T=32580 68120 0 0 $X=32500 $Y=67870
X135 28 M2_M1_CDNS_3 $T=33670 6150 0 90 $X=33420 $Y=6070
X136 26 M2_M1_CDNS_3 $T=34970 65150 0 0 $X=34890 $Y=64900
X137 19 M2_M1_CDNS_3 $T=34970 72470 0 0 $X=34890 $Y=72220
X138 10 M2_M1_CDNS_3 $T=37620 30320 0 0 $X=37540 $Y=30070
X139 33 M2_M1_CDNS_3 $T=40360 10220 0 90 $X=40110 $Y=10140
X140 33 M2_M1_CDNS_3 $T=40340 24940 0 0 $X=40260 $Y=24690
X141 33 M2_M1_CDNS_3 $T=40370 17590 0 0 $X=40290 $Y=17340
X142 12 M2_M1_CDNS_3 $T=40600 13810 0 0 $X=40520 $Y=13560
X143 32 M2_M1_CDNS_3 $T=40710 21060 0 0 $X=40630 $Y=20810
X144 15 M2_M1_CDNS_3 $T=46890 13630 0 0 $X=46810 $Y=13380
X145 15 M2_M1_CDNS_3 $T=46900 20740 0 0 $X=46820 $Y=20490
X146 15 M2_M1_CDNS_3 $T=46910 28080 0 0 $X=46830 $Y=27830
X147 33 M2_M1_CDNS_3 $T=47620 54480 0 90 $X=47370 $Y=54400
X148 33 M2_M1_CDNS_3 $T=47800 38230 0 90 $X=47550 $Y=38150
X149 33 M2_M1_CDNS_3 $T=47870 10240 0 0 $X=47790 $Y=9990
X150 33 M2_M1_CDNS_3 $T=47980 9490 0 180 $X=47900 $Y=9240
X151 33 M2_M1_CDNS_3 $T=48260 51950 0 90 $X=48010 $Y=51870
X152 33 M2_M1_CDNS_3 $T=48260 45130 0 0 $X=48180 $Y=44880
X153 33 M2_M1_CDNS_3 $T=48690 16910 0 0 $X=48610 $Y=16660
X154 33 M2_M1_CDNS_3 $T=48860 24230 0 0 $X=48780 $Y=23980
X155 33 M2_M1_CDNS_3 $T=48880 2280 0 0 $X=48800 $Y=2030
X156 1 M2_M1_CDNS_3 $T=49180 4060 0 0 $X=49100 $Y=3810
X157 1 M2_M1_CDNS_3 $T=49180 11470 0 0 $X=49100 $Y=11220
X158 1 M2_M1_CDNS_3 $T=49180 18800 0 0 $X=49100 $Y=18550
X159 1 M2_M1_CDNS_3 $T=49180 26120 0 0 $X=49100 $Y=25870
X160 1 M2_M1_CDNS_3 $T=49180 33430 0 0 $X=49100 $Y=33180
X161 1 M2_M1_CDNS_3 $T=49180 40820 0 0 $X=49100 $Y=40570
X162 1 M2_M1_CDNS_3 $T=49180 48070 0 0 $X=49100 $Y=47820
X163 1 M2_M1_CDNS_3 $T=49180 54710 0 0 $X=49100 $Y=54460
X164 13 M2_M1_CDNS_3 $T=50910 13780 0 0 $X=50830 $Y=13530
X165 17 M2_M1_CDNS_3 $T=58670 9650 0 90 $X=58420 $Y=9570
X166 17 M2_M1_CDNS_3 $T=58670 12550 0 90 $X=58420 $Y=12470
X167 17 M2_M1_CDNS_3 $T=58670 16970 0 90 $X=58420 $Y=16890
X168 17 M2_M1_CDNS_3 $T=58670 19870 0 90 $X=58420 $Y=19790
X169 17 M2_M1_CDNS_3 $T=58670 24290 0 90 $X=58420 $Y=24210
X170 17 M2_M1_CDNS_3 $T=58670 27190 0 90 $X=58420 $Y=27110
X171 17 M2_M1_CDNS_3 $T=58670 31610 0 90 $X=58420 $Y=31530
X172 17 M2_M1_CDNS_3 $T=58670 38930 0 90 $X=58420 $Y=38850
X173 17 M2_M1_CDNS_3 $T=58670 46250 0 90 $X=58420 $Y=46170
X174 17 M2_M1_CDNS_3 $T=58670 53570 0 90 $X=58420 $Y=53490
X175 14 M2_M1_CDNS_3 $T=59660 13790 0 0 $X=59580 $Y=13540
X176 30 M2_M1_CDNS_3 $T=59660 21120 0 0 $X=59580 $Y=20870
X177 28 M2_M1_CDNS_3 $T=59660 28470 0 0 $X=59580 $Y=28220
X178 18 M5_M4_CDNS_4 $T=1480 56760 0 0 $X=1400 $Y=56510
X179 19 M5_M4_CDNS_4 $T=2350 44590 0 90 $X=2100 $Y=44510
X180 20 M5_M4_CDNS_4 $T=3900 48300 0 90 $X=3650 $Y=48220
X181 21 M5_M4_CDNS_4 $T=3940 58210 0 90 $X=3690 $Y=58130
X182 18 M5_M4_CDNS_4 $T=4250 65060 0 180 $X=4170 $Y=64810
X183 21 M5_M4_CDNS_4 $T=4250 72470 0 0 $X=4170 $Y=72220
X184 22 M5_M4_CDNS_4 $T=6840 58120 0 90 $X=6590 $Y=58040
X185 23 M5_M4_CDNS_4 $T=11380 56560 0 90 $X=11130 $Y=56480
X186 23 M5_M4_CDNS_4 $T=14490 65150 0 0 $X=14410 $Y=64900
X187 22 M5_M4_CDNS_4 $T=14490 72480 0 0 $X=14410 $Y=72230
X188 24 M5_M4_CDNS_4 $T=20420 56560 0 90 $X=20170 $Y=56480
X189 24 M5_M4_CDNS_4 $T=24730 65150 0 0 $X=24650 $Y=64900
X190 20 M5_M4_CDNS_4 $T=24730 72470 0 0 $X=24650 $Y=72220
X191 25 M5_M4_CDNS_4 $T=27620 26990 0 0 $X=27540 $Y=26740
X192 26 M5_M4_CDNS_4 $T=29230 56560 0 90 $X=28980 $Y=56480
X193 25 M5_M4_CDNS_4 $T=32380 35710 0 90 $X=32130 $Y=35630
X194 27 M5_M4_CDNS_4 $T=32470 34080 0 90 $X=32220 $Y=34000
X195 27 M5_M4_CDNS_4 $T=33360 32510 0 90 $X=33110 $Y=32430
X196 28 M5_M4_CDNS_4 $T=33670 6150 0 90 $X=33420 $Y=6070
X197 34 M5_M4_CDNS_4 $T=33880 28620 0 0 $X=33800 $Y=28370
X198 29 M5_M4_CDNS_4 $T=34010 30140 0 0 $X=33930 $Y=29890
X199 11 M5_M4_CDNS_4 $T=34370 21060 0 0 $X=34290 $Y=20810
X200 26 M5_M4_CDNS_4 $T=34970 65150 0 0 $X=34890 $Y=64900
X201 19 M5_M4_CDNS_4 $T=34970 72470 0 0 $X=34890 $Y=72220
X202 29 M5_M4_CDNS_4 $T=35130 53970 0 0 $X=35050 $Y=53720
X203 31 M5_M4_CDNS_4 $T=36160 20250 0 0 $X=36080 $Y=20000
X204 35 M5_M4_CDNS_4 $T=36500 13950 0 0 $X=36420 $Y=13700
X205 36 M5_M4_CDNS_4 $T=37400 32460 0 0 $X=37320 $Y=32210
X206 8 M5_M4_CDNS_4 $T=37820 20120 0 0 $X=37740 $Y=19870
X207 30 M5_M4_CDNS_4 $T=38220 15840 0 0 $X=38140 $Y=15590
X208 28 M5_M4_CDNS_4 $T=38250 22590 0 0 $X=38170 $Y=22340
X209 31 M5_M4_CDNS_4 $T=38270 21170 0 0 $X=38190 $Y=20920
X210 35 M5_M4_CDNS_4 $T=40460 17040 0 90 $X=40210 $Y=16960
X211 8 M5_M4_CDNS_4 $T=40660 20120 0 90 $X=40410 $Y=20040
X212 37 M5_M4_CDNS_4 $T=40730 9730 0 90 $X=40480 $Y=9650
X213 9 M5_M4_CDNS_4 $T=40560 26320 0 0 $X=40480 $Y=26070
X214 36 M5_M4_CDNS_4 $T=42630 35130 0 90 $X=42380 $Y=35050
X215 14 M5_M4_CDNS_4 $T=47280 7640 0 90 $X=47030 $Y=7560
X216 30 M5_M4_CDNS_4 $T=47850 15290 0 0 $X=47770 $Y=15040
X217 28 M5_M4_CDNS_4 $T=47850 23870 0 0 $X=47770 $Y=23620
X218 15 M5_M4_CDNS_4 $T=47890 45870 0 0 $X=47810 $Y=45620
X219 33 M5_M4_CDNS_4 $T=47980 9490 0 180 $X=47900 $Y=9240
X220 33 M5_M4_CDNS_4 $T=48880 2280 0 0 $X=48800 $Y=2030
X221 15 M5_M4_CDNS_4 $T=50250 45640 0 90 $X=50000 $Y=45560
X222 14 M5_M4_CDNS_4 $T=59660 13790 0 0 $X=59580 $Y=13540
X223 30 M5_M4_CDNS_4 $T=59660 21120 0 0 $X=59580 $Y=20870
X224 28 M5_M4_CDNS_4 $T=59660 28470 0 0 $X=59580 $Y=28220
X225 18 M4_M3_CDNS_5 $T=1480 56760 0 0 $X=1400 $Y=56510
X226 19 M4_M3_CDNS_5 $T=2350 44590 0 90 $X=2100 $Y=44510
X227 20 M4_M3_CDNS_5 $T=3900 48300 0 90 $X=3650 $Y=48220
X228 21 M4_M3_CDNS_5 $T=3940 58210 0 90 $X=3690 $Y=58130
X229 18 M4_M3_CDNS_5 $T=4250 65060 0 180 $X=4170 $Y=64810
X230 21 M4_M3_CDNS_5 $T=4250 72470 0 0 $X=4170 $Y=72220
X231 22 M4_M3_CDNS_5 $T=6840 58120 0 90 $X=6590 $Y=58040
X232 23 M4_M3_CDNS_5 $T=11380 56560 0 90 $X=11130 $Y=56480
X233 23 M4_M3_CDNS_5 $T=14490 65150 0 0 $X=14410 $Y=64900
X234 22 M4_M3_CDNS_5 $T=14490 72480 0 0 $X=14410 $Y=72230
X235 24 M4_M3_CDNS_5 $T=20420 56560 0 90 $X=20170 $Y=56480
X236 24 M4_M3_CDNS_5 $T=24730 65150 0 0 $X=24650 $Y=64900
X237 20 M4_M3_CDNS_5 $T=24730 72470 0 0 $X=24650 $Y=72220
X238 25 M4_M3_CDNS_5 $T=27620 26990 0 0 $X=27540 $Y=26740
X239 26 M4_M3_CDNS_5 $T=29230 56560 0 90 $X=28980 $Y=56480
X240 27 M4_M3_CDNS_5 $T=32470 34080 0 90 $X=32220 $Y=34000
X241 28 M4_M3_CDNS_5 $T=33670 6150 0 90 $X=33420 $Y=6070
X242 26 M4_M3_CDNS_5 $T=34970 65150 0 0 $X=34890 $Y=64900
X243 19 M4_M3_CDNS_5 $T=34970 72470 0 0 $X=34890 $Y=72220
X244 29 M4_M3_CDNS_5 $T=35130 53970 0 0 $X=35050 $Y=53720
X245 30 M4_M3_CDNS_5 $T=38220 15840 0 0 $X=38140 $Y=15590
X246 28 M4_M3_CDNS_5 $T=38250 22590 0 0 $X=38170 $Y=22340
X247 31 M4_M3_CDNS_5 $T=38270 21170 0 0 $X=38190 $Y=20920
X248 14 M4_M3_CDNS_5 $T=47280 7640 0 90 $X=47030 $Y=7560
X249 30 M4_M3_CDNS_5 $T=47850 15290 0 0 $X=47770 $Y=15040
X250 28 M4_M3_CDNS_5 $T=47850 23870 0 0 $X=47770 $Y=23620
X251 33 M4_M3_CDNS_5 $T=47980 9490 0 180 $X=47900 $Y=9240
X252 33 M4_M3_CDNS_5 $T=48880 2280 0 0 $X=48800 $Y=2030
X253 15 M4_M3_CDNS_5 $T=50250 45640 0 90 $X=50000 $Y=45560
X254 14 M4_M3_CDNS_5 $T=59660 13790 0 0 $X=59580 $Y=13540
X255 30 M4_M3_CDNS_5 $T=59660 21120 0 0 $X=59580 $Y=20870
X256 28 M4_M3_CDNS_5 $T=59660 28470 0 0 $X=59580 $Y=28220
X257 33 M1_PO_CDNS_6 $T=1860 60810 0 0 $X=1760 $Y=60560
X258 33 M1_PO_CDNS_6 $T=1870 68120 0 0 $X=1770 $Y=67870
X259 19 M1_PO_CDNS_6 $T=2350 44590 0 90 $X=2100 $Y=44490
X260 20 M1_PO_CDNS_6 $T=3900 48300 0 90 $X=3650 $Y=48200
X261 21 M1_PO_CDNS_6 $T=3940 58210 0 90 $X=3690 $Y=58110
X262 22 M1_PO_CDNS_6 $T=6840 58120 0 90 $X=6590 $Y=58020
X263 33 M1_PO_CDNS_6 $T=12100 60800 0 0 $X=12000 $Y=60550
X264 33 M1_PO_CDNS_6 $T=12100 68120 0 0 $X=12000 $Y=67870
X265 33 M1_PO_CDNS_6 $T=22340 68120 0 0 $X=22240 $Y=67870
X266 33 M1_PO_CDNS_6 $T=22350 60800 0 0 $X=22250 $Y=60550
X267 33 M1_PO_CDNS_6 $T=32580 60800 0 0 $X=32480 $Y=60550
X268 33 M1_PO_CDNS_6 $T=32580 68120 0 0 $X=32480 $Y=67870
X269 28 M1_PO_CDNS_6 $T=33670 6150 0 90 $X=33420 $Y=6050
X270 33 M1_PO_CDNS_6 $T=40360 10220 0 90 $X=40110 $Y=10120
X271 33 M1_PO_CDNS_6 $T=40340 24940 0 0 $X=40240 $Y=24690
X272 33 M1_PO_CDNS_6 $T=40370 17590 0 0 $X=40270 $Y=17340
X273 15 M1_PO_CDNS_6 $T=46890 13630 0 0 $X=46790 $Y=13380
X274 15 M1_PO_CDNS_6 $T=46900 20740 0 0 $X=46800 $Y=20490
X275 15 M1_PO_CDNS_6 $T=46910 28080 0 0 $X=46810 $Y=27830
X276 33 M1_PO_CDNS_6 $T=47620 54480 0 90 $X=47370 $Y=54380
X277 33 M1_PO_CDNS_6 $T=47800 38230 0 90 $X=47550 $Y=38130
X278 33 M1_PO_CDNS_6 $T=47870 10240 0 0 $X=47770 $Y=9990
X279 33 M1_PO_CDNS_6 $T=47980 9490 0 180 $X=47880 $Y=9240
X280 33 M1_PO_CDNS_6 $T=48260 51950 0 90 $X=48010 $Y=51850
X281 33 M1_PO_CDNS_6 $T=48260 45130 0 0 $X=48160 $Y=44880
X282 33 M1_PO_CDNS_6 $T=48690 16910 0 0 $X=48590 $Y=16660
X283 33 M1_PO_CDNS_6 $T=48860 24230 0 0 $X=48760 $Y=23980
X284 33 M1_PO_CDNS_6 $T=48880 2280 0 0 $X=48780 $Y=2030
X285 3 M3_M2_CDNS_7 $T=15150 34320 0 0 $X=15070 $Y=34070
X286 5 M3_M2_CDNS_7 $T=30360 48950 0 0 $X=30280 $Y=48700
X287 6 M3_M2_CDNS_7 $T=30540 30290 0 90 $X=30290 $Y=30210
X288 7 M3_M2_CDNS_7 $T=30920 28440 0 90 $X=30670 $Y=28360
X289 7 M3_M2_CDNS_7 $T=30920 23090 0 0 $X=30840 $Y=22840
X290 6 M3_M2_CDNS_7 $T=30960 32190 0 0 $X=30880 $Y=31940
X291 8 M3_M2_CDNS_7 $T=34240 15510 0 0 $X=34160 $Y=15260
X292 9 M3_M2_CDNS_7 $T=36070 26280 0 0 $X=35990 $Y=26030
X293 6 M3_M2_CDNS_7 $T=36600 41550 0 0 $X=36520 $Y=41300
X294 11 M3_M2_CDNS_7 $T=37800 29000 0 0 $X=37720 $Y=28750
X295 12 M3_M2_CDNS_7 $T=40600 12040 0 0 $X=40520 $Y=11790
X296 13 M3_M2_CDNS_7 $T=41660 8130 0 0 $X=41580 $Y=7880
X297 14 M3_M2_CDNS_7 $T=43120 8620 0 0 $X=43040 $Y=8370
X298 15 M3_M2_CDNS_7 $T=45720 13840 0 0 $X=45640 $Y=13590
X299 15 M3_M2_CDNS_7 $T=47400 30300 0 0 $X=47320 $Y=30050
X300 16 M3_M2_CDNS_7 $T=50830 40760 0 90 $X=50580 $Y=40680
X301 17 M3_M2_CDNS_7 $T=58260 1650 0 0 $X=58180 $Y=1400
X302 32 M2_M1_CDNS_8 $T=13960 1790 0 90 $X=13830 $Y=1710
X303 3 M2_M1_CDNS_8 $T=26670 45180 0 0 $X=26590 $Y=45050
X304 36 M2_M1_CDNS_8 $T=27600 31220 0 0 $X=27520 $Y=31090
X305 38 M2_M1_CDNS_8 $T=28050 6240 0 0 $X=27970 $Y=6110
X306 8 M2_M1_CDNS_8 $T=28100 13310 0 0 $X=28020 $Y=13180
X307 13 M2_M1_CDNS_8 $T=28110 10050 0 0 $X=28030 $Y=9920
X308 9 M2_M1_CDNS_8 $T=28410 16430 0 90 $X=28280 $Y=16350
X309 27 M2_M1_CDNS_8 $T=35470 34490 0 0 $X=35390 $Y=34360
X310 12 M2_M1_CDNS_8 $T=35820 2210 0 90 $X=35690 $Y=2130
X311 7 M2_M1_CDNS_8 $T=37240 38080 0 0 $X=37160 $Y=37950
X312 38 M2_M1_CDNS_8 $T=41060 27730 0 0 $X=40980 $Y=27600
X313 5 M2_M1_CDNS_8 $T=43080 53380 0 0 $X=43000 $Y=53250
X314 15 M2_M1_CDNS_8 $T=47420 36740 0 0 $X=47340 $Y=36610
X315 10 M2_M1_CDNS_8 $T=47770 37090 0 0 $X=47690 $Y=36960
X316 25 M2_M1_CDNS_8 $T=50960 49840 0 90 $X=50830 $Y=49760
X317 16 M2_M1_CDNS_8 $T=51290 41540 0 90 $X=51160 $Y=41460
X318 8 M2_M1_CDNS_8 $T=51280 20630 0 0 $X=51200 $Y=20500
X319 4 M2_M1_CDNS_8 $T=51290 35200 0 0 $X=51210 $Y=35070
X320 9 M2_M1_CDNS_8 $T=51300 27960 0 0 $X=51220 $Y=27830
X321 36 M2_M1_CDNS_8 $T=51300 57100 0 0 $X=51220 $Y=56970
X322 37 M2_M1_CDNS_8 $T=59660 8330 0 0 $X=59580 $Y=8200
X323 35 M2_M1_CDNS_8 $T=59660 15640 0 0 $X=59580 $Y=15510
X324 31 M2_M1_CDNS_8 $T=59660 22940 0 0 $X=59580 $Y=22810
X325 11 M2_M1_CDNS_8 $T=59660 30310 0 0 $X=59580 $Y=30180
X326 10 M2_M1_CDNS_8 $T=59660 37620 0 0 $X=59580 $Y=37490
X327 34 M2_M1_CDNS_8 $T=59660 44940 0 0 $X=59580 $Y=44810
X328 29 M2_M1_CDNS_8 $T=59660 52270 0 0 $X=59580 $Y=52140
X329 33 M3_M2_CDNS_9 $T=1860 60810 0 0 $X=1780 $Y=60560
X330 33 M3_M2_CDNS_9 $T=1870 68120 0 0 $X=1790 $Y=67870
X331 33 M3_M2_CDNS_9 $T=12100 60800 0 0 $X=12020 $Y=60550
X332 33 M3_M2_CDNS_9 $T=12100 68120 0 0 $X=12020 $Y=67870
X333 33 M3_M2_CDNS_9 $T=22340 68120 0 0 $X=22260 $Y=67870
X334 33 M3_M2_CDNS_9 $T=22350 60800 0 0 $X=22270 $Y=60550
X335 39 M3_M2_CDNS_9 $T=22980 34240 0 0 $X=22900 $Y=33990
X336 16 M3_M2_CDNS_9 $T=28400 24370 0 0 $X=28320 $Y=24120
X337 40 M3_M2_CDNS_9 $T=32190 56290 0 0 $X=32110 $Y=56040
X338 33 M3_M2_CDNS_9 $T=32580 60800 0 0 $X=32500 $Y=60550
X339 33 M3_M2_CDNS_9 $T=32580 68120 0 0 $X=32500 $Y=67870
X340 33 M3_M2_CDNS_9 $T=40360 10220 0 90 $X=40110 $Y=10140
X341 33 M3_M2_CDNS_9 $T=40340 24940 0 0 $X=40260 $Y=24690
X342 33 M3_M2_CDNS_9 $T=40370 17590 0 0 $X=40290 $Y=17340
X343 10 M3_M2_CDNS_9 $T=45710 34580 0 0 $X=45630 $Y=34330
X344 33 M3_M2_CDNS_9 $T=47620 54480 0 90 $X=47370 $Y=54400
X345 33 M3_M2_CDNS_9 $T=47800 38230 0 90 $X=47550 $Y=38150
X346 33 M3_M2_CDNS_9 $T=47870 10240 0 0 $X=47790 $Y=9990
X347 33 M3_M2_CDNS_9 $T=48260 51950 0 90 $X=48010 $Y=51870
X348 33 M3_M2_CDNS_9 $T=48260 45130 0 0 $X=48180 $Y=44880
X349 33 M3_M2_CDNS_9 $T=48690 16910 0 0 $X=48610 $Y=16660
X350 33 M3_M2_CDNS_9 $T=48860 24230 0 0 $X=48780 $Y=23980
X351 30 M3_M2_CDNS_10 $T=14040 560 0 0 $X=13960 $Y=430
X352 32 M3_M2_CDNS_10 $T=22250 3160 0 0 $X=22170 $Y=3030
X353 30 M3_M2_CDNS_10 $T=23920 6540 0 0 $X=23840 $Y=6410
X354 40 M3_M2_CDNS_10 $T=25520 48970 0 0 $X=25440 $Y=48840
X355 7 M3_M2_CDNS_10 $T=27740 16660 0 0 $X=27660 $Y=16530
X356 6 M3_M2_CDNS_10 $T=28010 24010 0 0 $X=27930 $Y=23880
X357 36 M3_M2_CDNS_10 $T=31460 30680 0 90 $X=31330 $Y=30600
X358 40 M3_M2_CDNS_10 $T=32190 54030 0 0 $X=32110 $Y=53900
X359 27 M3_M2_CDNS_10 $T=36910 32510 0 0 $X=36830 $Y=32380
X360 27 M3_M2_CDNS_10 $T=37470 13030 0 0 $X=37390 $Y=12900
X361 38 M3_M2_CDNS_10 $T=37590 8380 0 90 $X=37460 $Y=8300
X362 38 M3_M2_CDNS_10 $T=38080 28430 0 0 $X=38000 $Y=28300
X363 10 M3_M2_CDNS_10 $T=39590 33870 0 0 $X=39510 $Y=33740
X364 25 M3_M2_CDNS_10 $T=40110 35670 0 90 $X=39980 $Y=35590
X365 4 M3_M2_CDNS_10 $T=42020 34330 0 0 $X=41940 $Y=34200
X366 34 M3_M2_CDNS_10 $T=45640 37660 0 0 $X=45560 $Y=37530
X367 33 M3_M2_CDNS_10 $T=47780 30450 0 0 $X=47700 $Y=30320
X368 33 M3_M2_CDNS_10 $T=47810 35930 0 0 $X=47730 $Y=35800
X369 8 M3_M2_CDNS_10 $T=48170 20860 0 0 $X=48090 $Y=20730
X370 9 M3_M2_CDNS_10 $T=48180 28260 0 0 $X=48100 $Y=28130
X371 15 M3_M2_CDNS_10 $T=48350 54060 0 0 $X=48270 $Y=53930
X372 35 M3_M2_CDNS_10 $T=48430 15830 0 0 $X=48350 $Y=15700
X373 36 M3_M2_CDNS_10 $T=49580 57720 0 90 $X=49450 $Y=57640
X374 37 M3_M2_CDNS_10 $T=50600 8490 0 0 $X=50520 $Y=8360
X375 25 M4_M3_CDNS_11 $T=32380 35710 0 90 $X=32130 $Y=35630
X376 27 M4_M3_CDNS_11 $T=33360 32510 0 90 $X=33110 $Y=32430
X377 34 M4_M3_CDNS_11 $T=33880 28620 0 0 $X=33800 $Y=28370
X378 29 M4_M3_CDNS_11 $T=34010 30140 0 0 $X=33930 $Y=29890
X379 11 M4_M3_CDNS_11 $T=34370 21060 0 0 $X=34290 $Y=20810
X380 31 M4_M3_CDNS_11 $T=36160 20250 0 0 $X=36080 $Y=20000
X381 35 M4_M3_CDNS_11 $T=36500 13950 0 0 $X=36420 $Y=13700
X382 36 M4_M3_CDNS_11 $T=37400 32460 0 0 $X=37320 $Y=32210
X383 8 M4_M3_CDNS_11 $T=37820 20120 0 0 $X=37740 $Y=19870
X384 35 M4_M3_CDNS_11 $T=40460 17040 0 90 $X=40210 $Y=16960
X385 8 M4_M3_CDNS_11 $T=40660 20120 0 90 $X=40410 $Y=20040
X386 37 M4_M3_CDNS_11 $T=40730 9730 0 90 $X=40480 $Y=9650
X387 9 M4_M3_CDNS_11 $T=40560 26320 0 0 $X=40480 $Y=26070
X388 36 M4_M3_CDNS_11 $T=42630 35130 0 90 $X=42380 $Y=35050
X389 15 M4_M3_CDNS_11 $T=47890 45870 0 0 $X=47810 $Y=45620
X390 2 M4_M3_CDNS_12 $T=13710 9140 0 0 $X=13630 $Y=9010
X391 2 M4_M3_CDNS_12 $T=13710 17480 0 0 $X=13630 $Y=17350
X392 2 M4_M3_CDNS_12 $T=13710 19960 0 0 $X=13630 $Y=19830
X393 3 M4_M3_CDNS_12 $T=14090 21060 0 0 $X=14010 $Y=20930
X394 40 M4_M3_CDNS_12 $T=24590 43490 0 0 $X=24510 $Y=43360
X395 5 M4_M3_CDNS_12 $T=28000 27530 0 0 $X=27920 $Y=27400
X396 40 M4_M3_CDNS_12 $T=28120 30940 0 0 $X=28040 $Y=30810
X397 30 M4_M3_CDNS_12 $T=30320 6550 0 0 $X=30240 $Y=6420
X398 28 M4_M3_CDNS_12 $T=31030 8560 0 90 $X=30900 $Y=8480
X399 37 M4_M3_CDNS_12 $T=34270 8400 0 0 $X=34190 $Y=8270
X400 10 M4_M3_CDNS_12 $T=34570 23190 0 0 $X=34490 $Y=23060
X401 28 M4_M3_CDNS_12 $T=34690 12200 0 0 $X=34610 $Y=12070
X402 16 M4_M3_CDNS_12 $T=36100 30140 0 0 $X=36020 $Y=30010
X403 34 M4_M3_CDNS_12 $T=36540 37650 0 90 $X=36410 $Y=37570
X404 8 M4_M3_CDNS_12 $T=37250 15560 0 0 $X=37170 $Y=15430
X405 4 M4_M3_CDNS_12 $T=37310 22870 0 0 $X=37230 $Y=22740
X406 38 M4_M3_CDNS_12 $T=37550 19040 0 0 $X=37470 $Y=18910
X407 38 M4_M3_CDNS_12 $T=37670 21700 0 0 $X=37590 $Y=21570
X408 32 M4_M3_CDNS_12 $T=38370 9550 0 0 $X=38290 $Y=9420
X409 32 M4_M3_CDNS_12 $T=40710 21060 0 0 $X=40630 $Y=20930
X410 14 M4_M3_CDNS_12 $T=41120 2720 0 0 $X=41040 $Y=2590
X411 15 M4_M3_CDNS_12 $T=47400 30300 0 0 $X=47320 $Y=30170
X412 33 M4_M3_CDNS_12 $T=48170 14160 0 0 $X=48090 $Y=14030
X413 33 M4_M3_CDNS_12 $T=48170 17210 0 0 $X=48090 $Y=17080
X414 13 M4_M3_CDNS_12 $T=50910 13780 0 0 $X=50830 $Y=13650
X415 2 M2_M1_CDNS_13 $T=14700 34240 0 0 $X=14620 $Y=33990
X416 39 M2_M1_CDNS_13 $T=22980 34240 0 0 $X=22900 $Y=33990
X417 16 M2_M1_CDNS_13 $T=28400 24370 0 0 $X=28320 $Y=24120
X418 40 M2_M1_CDNS_13 $T=32190 56290 0 0 $X=32110 $Y=56040
X419 6 M2_M1_CDNS_13 $T=38820 45300 0 0 $X=38740 $Y=45050
X420 10 M2_M1_CDNS_13 $T=45710 34580 0 0 $X=45630 $Y=34330
X421 28 M5_M4_CDNS_14 $T=31030 6520 0 0 $X=30950 $Y=6390
X422 29 M5_M4_CDNS_14 $T=33450 34810 0 0 $X=33370 $Y=34680
X423 29 M5_M4_CDNS_14 $T=34490 38940 0 0 $X=34410 $Y=38810
X424 29 M5_M4_CDNS_14 $T=35140 50450 0 0 $X=35060 $Y=50320
X425 11 M5_M4_CDNS_14 $T=35270 23970 0 0 $X=35190 $Y=23840
X426 29 M5_M4_CDNS_14 $T=35630 42220 0 0 $X=35550 $Y=42090
X427 28 M5_M4_CDNS_14 $T=35740 16590 0 0 $X=35660 $Y=16460
X428 34 M5_M4_CDNS_14 $T=36550 34300 0 0 $X=36470 $Y=34170
X429 16 M5_M4_CDNS_14 $T=36920 33010 0 0 $X=36840 $Y=32880
X430 30 M5_M4_CDNS_14 $T=37650 13930 0 0 $X=37570 $Y=13800
X431 37 M5_M4_CDNS_14 $T=37800 9740 0 0 $X=37720 $Y=9610
X432 14 M5_M4_CDNS_14 $T=38000 8190 0 0 $X=37920 $Y=8060
X433 32 M5_M4_CDNS_14 $T=38690 18860 0 90 $X=38560 $Y=18780
X434 9 M5_M4_CDNS_14 $T=38750 26290 0 90 $X=38620 $Y=26210
X435 32 M5_M4_CDNS_14 $T=40200 18860 0 90 $X=40070 $Y=18780
X436 14 M5_M4_CDNS_14 $T=40300 8620 0 90 $X=40170 $Y=8540
X437 13 M5_M4_CDNS_14 $T=48360 8140 0 0 $X=48280 $Y=8010
X438 13 M5_M4_CDNS_14 $T=50330 8160 0 0 $X=50250 $Y=8030
X439 16 M5_M4_CDNS_14 $T=50340 37430 0 0 $X=50260 $Y=37300
X440 33 M1_PO_CDNS_15 $T=47780 31470 0 0 $X=47680 $Y=31220
X441 15 M1_PO_CDNS_16 $T=47950 48930 0 0 $X=47850 $Y=48810
X442 33 M2_M1_CDNS_17 $T=47780 31470 0 0 $X=47700 $Y=31220
X443 18 1 21 20 19 41 23 24 22 2
+ 26 39 3 40 27 7 6 5 92 93
+ 139 77 150 79 140 151 127 138 136 178
+ 154 179 168 111 114 174 112 75 121 110
+ 175 157 80 161 123 177 89 85 149 122 multiplier $T=1090 33260 0 0 $X=750 $Y=33040
X444 30 42 41 1 43 7 40 28 37 35
+ 11 10 34 29 5 6 3 31 27 2
+ 39 32 14 44 36 4 16 25 38 13
+ 8 9 12 45 193 203 202 239 309 208
+ 207 210 209 213 212 219 218 217 216 201
+ 200 205 204 195 194 197 196 199 198 10badder $T=-50390 53780 1 0 $X=-110 $Y=0
X445 41 15 1 33 18 46 318 315 683 316
+ 685 314 319 312 313 317 320 ph1p3_MSDFF $T=1140 62320 0 0 $X=1140 $Y=58560
X446 41 15 1 33 21 47 327 324 686 325
+ 688 323 328 321 322 326 329 ph1p3_MSDFF $T=1140 69640 0 0 $X=1140 $Y=65880
X447 41 15 1 33 23 48 336 333 689 334
+ 691 332 337 330 331 335 338 ph1p3_MSDFF $T=11380 62320 0 0 $X=11380 $Y=58560
X448 41 15 1 33 22 49 345 342 692 343
+ 694 341 346 339 340 344 347 ph1p3_MSDFF $T=11380 69640 0 0 $X=11380 $Y=65880
X449 41 15 1 33 24 50 354 351 695 352
+ 697 350 355 348 349 353 356 ph1p3_MSDFF $T=21620 62320 0 0 $X=21620 $Y=58560
X450 41 15 1 33 20 51 363 360 698 361
+ 700 359 364 357 358 362 365 ph1p3_MSDFF $T=21620 69640 0 0 $X=21620 $Y=65880
X451 41 15 1 33 26 52 372 369 701 370
+ 703 368 373 366 367 371 374 ph1p3_MSDFF $T=31860 62320 0 0 $X=31860 $Y=58560
X452 41 15 1 33 19 53 381 378 704 379
+ 706 377 382 375 376 380 383 ph1p3_MSDFF $T=31860 69640 0 0 $X=31860 $Y=65880
X453 41 15 1 33 12 14 390 387 707 388
+ 709 386 391 384 385 389 392 ph1p3_MSDFF $T=37920 11080 0 0 $X=37920 $Y=7320
X454 41 15 1 33 32 30 399 396 710 397
+ 712 395 400 393 394 398 401 ph1p3_MSDFF $T=37920 18400 0 0 $X=37920 $Y=14640
X455 41 15 1 33 38 28 408 405 713 406
+ 715 404 409 402 403 407 410 ph1p3_MSDFF $T=37920 25720 0 0 $X=37920 $Y=21960
X456 41 15 1 33 54 17 417 414 716 415
+ 718 413 418 411 412 416 419 ph1p3_MSDFF $T=48160 3760 0 0 $X=48160 $Y=0
X457 41 15 1 33 13 37 426 423 719 424
+ 721 422 427 420 421 425 428 ph1p3_MSDFF $T=48160 11080 0 0 $X=48160 $Y=7320
X458 41 15 1 33 8 35 435 432 722 433
+ 724 431 436 429 430 434 437 ph1p3_MSDFF $T=48160 18400 0 0 $X=48160 $Y=14640
X459 41 15 1 33 9 31 444 441 725 442
+ 727 440 445 438 439 443 446 ph1p3_MSDFF $T=48160 25720 0 0 $X=48160 $Y=21960
X460 41 15 1 33 4 11 453 450 728 451
+ 730 449 454 447 448 452 455 ph1p3_MSDFF $T=48160 33040 0 0 $X=48160 $Y=29280
X461 41 15 1 33 16 10 462 459 731 460
+ 733 458 463 456 457 461 464 ph1p3_MSDFF $T=48160 40360 0 0 $X=48160 $Y=36600
X462 41 15 1 33 25 34 471 468 734 469
+ 736 467 472 465 466 470 473 ph1p3_MSDFF $T=48160 47680 0 0 $X=48160 $Y=43920
X463 41 15 1 33 36 29 480 477 737 478
+ 739 476 481 474 475 479 482 ph1p3_MSDFF $T=48160 55000 0 0 $X=48160 $Y=51240
X464 41 1 cellTmpl_CDNS_49 $T=47620 54900 1 0 $X=47500 $Y=51240
X465 17 37 41 1 55 56 483 484 740 741
+ 766 767 MUX_2to1___2X_ph2p2 $T=58160 11120 1 0 $X=58160 $Y=7320
X466 17 14 41 1 57 58 485 486 742 743
+ 768 769 MUX_2to1___2X_ph2p2 $T=58160 11080 0 0 $X=58160 $Y=11080
X467 17 35 41 1 59 60 487 488 744 745
+ 770 771 MUX_2to1___2X_ph2p2 $T=58160 18440 1 0 $X=58160 $Y=14640
X468 17 30 41 1 61 62 489 490 746 747
+ 772 773 MUX_2to1___2X_ph2p2 $T=58160 18400 0 0 $X=58160 $Y=18400
X469 17 31 41 1 63 64 491 492 748 749
+ 774 775 MUX_2to1___2X_ph2p2 $T=58160 25760 1 0 $X=58160 $Y=21960
X470 17 28 41 1 65 66 493 494 750 751
+ 776 777 MUX_2to1___2X_ph2p2 $T=58160 25720 0 0 $X=58160 $Y=25720
X471 17 11 41 1 67 68 495 496 752 753
+ 778 779 MUX_2to1___2X_ph2p2 $T=58160 33080 1 0 $X=58160 $Y=29280
X472 17 10 41 1 69 70 497 498 754 755
+ 780 781 MUX_2to1___2X_ph2p2 $T=58160 40400 1 0 $X=58160 $Y=36600
X473 17 34 41 1 71 72 499 500 756 757
+ 782 783 MUX_2to1___2X_ph2p2 $T=58160 47720 1 0 $X=58160 $Y=43920
X474 17 29 41 1 73 74 501 502 758 759
+ 784 785 MUX_2to1___2X_ph2p2 $T=58160 55040 1 0 $X=58160 $Y=51240
M0 315 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=59450 $dt=1
M1 318 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=64750 $dt=1
M2 324 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=66770 $dt=1
M3 327 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=1920 $Y=72070 $dt=1
M4 312 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3250 $Y=64780 $dt=1
M5 321 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=3250 $Y=72100 $dt=1
M6 313 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=59420 $dt=1
M7 322 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=66740 $dt=1
M8 314 15 18 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4430 $Y=64780 $dt=1
M9 323 15 21 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=4430 $Y=72100 $dt=1
M10 319 15 683 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=59660 $dt=1
M11 328 15 686 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=66980 $dt=1
M12 316 314 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5630 $Y=64690 $dt=1
M13 325 323 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=5630 $Y=72010 $dt=1
M14 683 46 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=59450 $dt=1
M15 686 47 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=66770 $dt=1
M16 316 315 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6870 $Y=64700 $dt=1
M17 325 324 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=6870 $Y=72020 $dt=1
M18 317 318 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=59420 $dt=1
M19 326 327 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=66740 $dt=1
M20 685 316 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8120 $Y=64750 $dt=1
M21 688 325 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=8120 $Y=72070 $dt=1
M22 319 318 316 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=59660 $dt=1
M23 328 327 325 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=66980 $dt=1
M24 320 318 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9450 $Y=64780 $dt=1
M25 329 327 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=9450 $Y=72100 $dt=1
M26 46 319 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=59450 $dt=1
M27 47 328 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=66770 $dt=1
M28 314 318 685 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=10630 $Y=64780 $dt=1
M29 323 327 688 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=10630 $Y=72100 $dt=1
M30 333 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=59450 $dt=1
M31 336 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=64750 $dt=1
M32 342 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=66770 $dt=1
M33 345 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=12160 $Y=72070 $dt=1
M34 330 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13490 $Y=64780 $dt=1
M35 339 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=13490 $Y=72100 $dt=1
M36 331 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=59420 $dt=1
M37 340 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=66740 $dt=1
M38 332 15 23 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=14670 $Y=64780 $dt=1
M39 341 15 22 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=14670 $Y=72100 $dt=1
M40 337 15 689 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=59660 $dt=1
M41 346 15 692 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=66980 $dt=1
M42 334 332 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=15870 $Y=64690 $dt=1
M43 343 341 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=15870 $Y=72010 $dt=1
M44 689 48 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=59450 $dt=1
M45 692 49 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=66770 $dt=1
M46 334 333 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17110 $Y=64700 $dt=1
M47 343 342 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=17110 $Y=72020 $dt=1
M48 335 336 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=59420 $dt=1
M49 344 345 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=66740 $dt=1
M50 691 334 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18360 $Y=64750 $dt=1
M51 694 343 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=18360 $Y=72070 $dt=1
M52 337 336 334 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=59660 $dt=1
M53 346 345 343 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=66980 $dt=1
M54 338 336 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=19690 $Y=64780 $dt=1
M55 347 345 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=19690 $Y=72100 $dt=1
M56 48 337 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=59450 $dt=1
M57 49 346 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=66770 $dt=1
M58 332 336 691 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=20870 $Y=64780 $dt=1
M59 341 345 694 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=20870 $Y=72100 $dt=1
M60 351 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=59450 $dt=1
M61 354 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=64750 $dt=1
M62 360 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=66770 $dt=1
M63 363 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=22400 $Y=72070 $dt=1
M64 348 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=23730 $Y=64780 $dt=1
M65 357 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=23730 $Y=72100 $dt=1
M66 349 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=59420 $dt=1
M67 358 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=66740 $dt=1
M68 350 15 24 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=24910 $Y=64780 $dt=1
M69 359 15 20 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=24910 $Y=72100 $dt=1
M70 355 15 695 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=59660 $dt=1
M71 364 15 698 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=66980 $dt=1
M72 352 350 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26110 $Y=64690 $dt=1
M73 361 359 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=26110 $Y=72010 $dt=1
M74 695 50 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=59450 $dt=1
M75 698 51 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=66770 $dt=1
M76 352 351 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27350 $Y=64700 $dt=1
M77 361 360 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=27350 $Y=72020 $dt=1
M78 353 354 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=59420 $dt=1
M79 362 363 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=66740 $dt=1
M80 697 352 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28600 $Y=64750 $dt=1
M81 700 361 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=28600 $Y=72070 $dt=1
M82 355 354 352 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=59660 $dt=1
M83 364 363 361 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=66980 $dt=1
M84 356 354 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=29930 $Y=64780 $dt=1
M85 365 363 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=29930 $Y=72100 $dt=1
M86 50 355 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=59450 $dt=1
M87 51 364 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=66770 $dt=1
M88 350 354 697 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31110 $Y=64780 $dt=1
M89 359 363 700 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=31110 $Y=72100 $dt=1
M90 369 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=59450 $dt=1
M91 372 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=64750 $dt=1
M92 378 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=66770 $dt=1
M93 381 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=32640 $Y=72070 $dt=1
M94 366 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=33970 $Y=64780 $dt=1
M95 375 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=33970 $Y=72100 $dt=1
M96 367 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=59420 $dt=1
M97 376 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=66740 $dt=1
M98 368 15 26 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35150 $Y=64780 $dt=1
M99 377 15 19 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=35150 $Y=72100 $dt=1
M100 373 15 701 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=59660 $dt=1
M101 382 15 704 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=66980 $dt=1
M102 370 368 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36350 $Y=64690 $dt=1
M103 379 377 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=36350 $Y=72010 $dt=1
M104 701 52 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=37440 $Y=59450 $dt=1
M105 704 53 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=37440 $Y=66770 $dt=1
M106 370 369 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37590 $Y=64700 $dt=1
M107 379 378 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=37590 $Y=72020 $dt=1
M108 387 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=8210 $dt=1
M109 390 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=13510 $dt=1
M110 396 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=15530 $dt=1
M111 399 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=20830 $dt=1
M112 405 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=22850 $dt=1
M113 408 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=28150 $dt=1
M114 371 372 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=38770 $Y=59420 $dt=1
M115 380 381 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=38770 $Y=66740 $dt=1
M116 703 370 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=38840 $Y=64750 $dt=1
M117 706 379 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=38840 $Y=72070 $dt=1
M118 373 372 370 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=39950 $Y=59660 $dt=1
M119 382 381 379 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=39950 $Y=66980 $dt=1
M120 384 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=13540 $dt=1
M121 393 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=20860 $dt=1
M122 402 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=40030 $Y=28180 $dt=1
M123 374 372 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40170 $Y=64780 $dt=1
M124 383 381 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=40170 $Y=72100 $dt=1
M125 385 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=41030 $Y=8180 $dt=1
M126 394 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=15500 $dt=1
M127 403 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=22820 $dt=1
M128 386 15 12 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=13540 $dt=1
M129 395 15 32 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=20860 $dt=1
M130 404 15 38 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=41210 $Y=28180 $dt=1
M131 52 373 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=41240 $Y=59450 $dt=1
M132 53 382 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=41240 $Y=66770 $dt=1
M133 368 372 703 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41350 $Y=64780 $dt=1
M134 377 381 706 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=41350 $Y=72100 $dt=1
M135 391 15 707 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=42210 $Y=8420 $dt=1
M136 400 15 710 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=15740 $dt=1
M137 409 15 713 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=23060 $dt=1
M138 388 386 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=13450 $dt=1
M139 397 395 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=20770 $dt=1
M140 406 404 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42410 $Y=28090 $dt=1
M141 707 14 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=43500 $Y=8210 $dt=1
M142 710 30 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=15530 $dt=1
M143 713 28 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=22850 $dt=1
M144 388 387 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=13460 $dt=1
M145 397 396 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=20780 $dt=1
M146 406 405 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43650 $Y=28100 $dt=1
M147 389 390 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=44830 $Y=8180 $dt=1
M148 398 399 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=15500 $dt=1
M149 407 408 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=22820 $dt=1
M150 709 388 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=13510 $dt=1
M151 712 397 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=20830 $dt=1
M152 715 406 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=44900 $Y=28150 $dt=1
M153 391 390 388 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=46010 $Y=8420 $dt=1
M154 400 399 397 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=15740 $dt=1
M155 409 408 406 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=23060 $dt=1
M156 392 390 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=13540 $dt=1
M157 401 399 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=20860 $dt=1
M158 410 408 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=46230 $Y=28180 $dt=1
M159 14 391 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=47300 $Y=8210 $dt=1
M160 30 400 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=15530 $dt=1
M161 28 409 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=22850 $dt=1
M162 386 390 709 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=13540 $dt=1
M163 395 399 712 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=20860 $dt=1
M164 404 408 715 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=47410 $Y=28180 $dt=1
M165 414 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=890 $dt=1
M166 417 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=6190 $dt=1
M167 423 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=8210 $dt=1
M168 426 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=13510 $dt=1
M169 432 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=15530 $dt=1
M170 435 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=20830 $dt=1
M171 441 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=22850 $dt=1
M172 444 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=28150 $dt=1
M173 450 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=30170 $dt=1
M174 453 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=35470 $dt=1
M175 459 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=37490 $dt=1
M176 462 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=42790 $dt=1
M177 468 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=44810 $dt=1
M178 471 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=50110 $dt=1
M179 477 33 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=52130 $dt=1
M180 480 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=57430 $dt=1
M181 411 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=6220 $dt=1
M182 420 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=13540 $dt=1
M183 429 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=20860 $dt=1
M184 438 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=28180 $dt=1
M185 447 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=35500 $dt=1
M186 456 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=42820 $dt=1
M187 465 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=50140 $dt=1
M188 474 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=50270 $Y=57460 $dt=1
M189 412 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=51270 $Y=860 $dt=1
M190 421 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=8180 $dt=1
M191 430 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=15500 $dt=1
M192 439 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=22820 $dt=1
M193 448 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=30140 $dt=1
M194 457 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=37460 $dt=1
M195 466 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=44780 $dt=1
M196 475 15 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=52100 $dt=1
M197 413 15 54 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=6220 $dt=1
M198 422 15 13 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=13540 $dt=1
M199 431 15 8 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=20860 $dt=1
M200 440 15 9 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=28180 $dt=1
M201 449 15 4 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=35500 $dt=1
M202 458 15 16 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=42820 $dt=1
M203 467 15 25 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=50140 $dt=1
M204 476 15 36 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=51450 $Y=57460 $dt=1
M205 418 15 716 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=52450 $Y=1100 $dt=1
M206 427 15 719 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=8420 $dt=1
M207 436 15 722 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=15740 $dt=1
M208 445 15 725 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=23060 $dt=1
M209 454 15 728 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=30380 $dt=1
M210 463 15 731 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=37700 $dt=1
M211 472 15 734 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=45020 $dt=1
M212 481 15 737 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=52340 $dt=1
M213 415 413 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=6130 $dt=1
M214 424 422 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=13450 $dt=1
M215 433 431 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=20770 $dt=1
M216 442 440 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=28090 $dt=1
M217 451 449 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=35410 $dt=1
M218 460 458 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=42730 $dt=1
M219 469 467 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=50050 $dt=1
M220 478 476 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=52650 $Y=57370 $dt=1
M221 716 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=53740 $Y=890 $dt=1
M222 719 37 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=8210 $dt=1
M223 722 35 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=15530 $dt=1
M224 725 31 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=22850 $dt=1
M225 728 11 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=30170 $dt=1
M226 731 10 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=37490 $dt=1
M227 734 34 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=44810 $dt=1
M228 737 29 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=52130 $dt=1
M229 415 414 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=6140 $dt=1
M230 424 423 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=13460 $dt=1
M231 433 432 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=20780 $dt=1
M232 442 441 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=28100 $dt=1
M233 451 450 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=35420 $dt=1
M234 460 459 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=42740 $dt=1
M235 469 468 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=50060 $dt=1
M236 478 477 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=53890 $Y=57380 $dt=1
M237 416 417 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=55070 $Y=860 $dt=1
M238 425 426 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=8180 $dt=1
M239 434 435 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=15500 $dt=1
M240 443 444 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=22820 $dt=1
M241 452 453 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=30140 $dt=1
M242 461 462 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=37460 $dt=1
M243 470 471 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=44780 $dt=1
M244 479 480 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=52100 $dt=1
M245 718 415 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=6190 $dt=1
M246 721 424 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=13510 $dt=1
M247 724 433 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=20830 $dt=1
M248 727 442 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=28150 $dt=1
M249 730 451 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=35470 $dt=1
M250 733 460 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=42790 $dt=1
M251 736 469 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=50110 $dt=1
M252 739 478 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=55140 $Y=57430 $dt=1
M253 418 417 415 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=56250 $Y=1100 $dt=1
M254 427 426 424 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=8420 $dt=1
M255 436 435 433 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=15740 $dt=1
M256 445 444 442 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=23060 $dt=1
M257 454 453 451 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=30380 $dt=1
M258 463 462 460 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=37700 $dt=1
M259 472 471 469 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=45020 $dt=1
M260 481 480 478 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=52340 $dt=1
M261 419 417 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=6220 $dt=1
M262 428 426 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=13540 $dt=1
M263 437 435 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=20860 $dt=1
M264 446 444 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=28180 $dt=1
M265 455 453 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=35500 $dt=1
M266 464 462 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=42820 $dt=1
M267 473 471 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=50140 $dt=1
M268 482 480 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=56470 $Y=57460 $dt=1
M269 17 418 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=57540 $Y=890 $dt=1
M270 37 427 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=8210 $dt=1
M271 35 436 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=15530 $dt=1
M272 31 445 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=22850 $dt=1
M273 11 454 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=30170 $dt=1
M274 10 463 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=37490 $dt=1
M275 34 472 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=44810 $dt=1
M276 29 481 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=52130 $dt=1
M277 413 417 718 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=6220 $dt=1
M278 422 426 721 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=13540 $dt=1
M279 431 435 724 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=20860 $dt=1
M280 440 444 727 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=28180 $dt=1
M281 449 453 730 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=35500 $dt=1
M282 458 462 733 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=42820 $dt=1
M283 467 471 736 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=50140 $dt=1
M284 476 480 739 41 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=57650 $Y=57460 $dt=1
M285 483 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=8270 $dt=1
M286 485 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=13450 $dt=1
M287 487 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=15590 $dt=1
M288 489 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=20770 $dt=1
M289 491 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=22910 $dt=1
M290 493 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=28090 $dt=1
M291 495 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=30230 $dt=1
M292 497 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=37550 $dt=1
M293 499 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=44870 $dt=1
M294 501 17 41 41 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=52190 $dt=1
M295 766 37 484 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=8060 $dt=1
M296 768 14 486 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=13180 $dt=1
M297 770 35 488 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=15380 $dt=1
M298 772 30 490 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=20500 $dt=1
M299 774 31 492 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=22700 $dt=1
M300 776 28 494 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=27820 $dt=1
M301 778 11 496 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=30020 $dt=1
M302 780 10 498 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=37340 $dt=1
M303 782 34 500 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=44660 $dt=1
M304 784 29 502 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=51980 $dt=1
M305 41 17 766 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=8060 $dt=1
M306 41 17 768 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=13180 $dt=1
M307 41 17 770 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=15380 $dt=1
M308 41 17 772 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=20500 $dt=1
M309 41 17 774 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=22700 $dt=1
M310 41 17 776 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=27820 $dt=1
M311 41 17 778 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=30020 $dt=1
M312 41 17 780 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=37340 $dt=1
M313 41 17 782 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=44660 $dt=1
M314 41 17 784 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=51980 $dt=1
M315 767 483 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=8130 $dt=1
M316 769 485 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=13110 $dt=1
M317 771 487 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=15450 $dt=1
M318 773 489 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=20430 $dt=1
M319 775 491 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=22770 $dt=1
M320 777 493 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=27750 $dt=1
M321 779 495 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=30090 $dt=1
M322 781 497 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=37410 $dt=1
M323 783 499 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=44730 $dt=1
M324 785 501 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=52050 $dt=1
M325 484 55 767 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=8130 $dt=1
M326 486 57 769 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=13110 $dt=1
M327 488 59 771 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=15450 $dt=1
M328 490 61 773 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=20430 $dt=1
M329 492 63 775 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=22770 $dt=1
M330 494 65 777 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=27750 $dt=1
M331 496 67 779 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=30090 $dt=1
M332 498 69 781 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=37410 $dt=1
M333 500 71 783 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=44730 $dt=1
M334 502 73 785 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=52050 $dt=1
M335 56 484 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=8120 $dt=1
M336 58 486 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=13120 $dt=1
M337 60 488 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=15440 $dt=1
M338 62 490 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=20440 $dt=1
M339 64 492 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=22760 $dt=1
M340 66 494 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=27760 $dt=1
M341 68 496 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=30080 $dt=1
M342 70 498 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=37400 $dt=1
M343 72 500 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=44720 $dt=1
M344 74 502 41 41 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=52040 $dt=1
.ends ph2p2_processing_element
