* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph1p3_DFF                                    *
* Netlisted  : Thu Nov  7 22:31:47 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_7                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_7 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 1 M1_PO_CDNS_6 $T=700 2040 0 90 $X=580 $Y=1940
X1 2 3 cellTmpl_CDNS_7 $T=120 140 0 0 $X=0 $Y=0
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=780 $Y=900 $dt=0
.ends INV_1X_small_layout

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_8                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_8 1 2 3 4
** N=4 EP=4 FDC=1
M0 2 3 1 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_9                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_9 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_11                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_11 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_6 $T=640 1830 0 90 $X=520 $Y=1730
X1 6 M1_PO_CDNS_6 $T=1940 640 0 0 $X=1840 $Y=520
X2 3 6 1 3 nmos1v_CDNS_8 $T=710 860 0 0 $X=290 $Y=660
X3 4 5 6 3 nmos1v_CDNS_8 $T=1890 860 0 0 $X=1470 $Y=660
X4 2 6 1 3 2 pmos1v_CDNS_9 $T=710 2460 0 0 $X=290 $Y=2260
X5 4 5 1 3 2 pmos1v_CDNS_11 $T=1890 2460 0 0 $X=1470 $Y=2260
.ends ph1p3_clk_part

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_DFF                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_DFF 4 11 6 10 9
** N=15 EP=5 FDC=26
X0 1 M3_M2_CDNS_1 $T=1220 2180 0 90 $X=970 $Y=2100
X1 2 M3_M2_CDNS_1 $T=3460 -2020 0 0 $X=3380 $Y=-2270
X2 3 M3_M2_CDNS_1 $T=4010 1790 0 0 $X=3930 $Y=1540
X3 1 M3_M2_CDNS_1 $T=5640 -1640 0 0 $X=5560 $Y=-1890
X4 1 M3_M2_CDNS_1 $T=7110 2180 0 90 $X=6860 $Y=2100
X5 2 M3_M2_CDNS_1 $T=7750 -1970 0 0 $X=7670 $Y=-2220
X6 3 M3_M2_CDNS_1 $T=8830 1770 0 0 $X=8750 $Y=1520
X7 1 M2_M1_CDNS_4 $T=1220 2180 0 90 $X=970 $Y=2100
X8 2 M2_M1_CDNS_4 $T=3460 -2020 0 0 $X=3380 $Y=-2270
X9 3 M2_M1_CDNS_4 $T=4010 1790 0 0 $X=3930 $Y=1540
X10 1 M2_M1_CDNS_4 $T=5640 -1640 0 0 $X=5560 $Y=-1890
X11 2 M2_M1_CDNS_4 $T=7750 -1970 0 0 $X=7670 $Y=-2220
X12 3 M2_M1_CDNS_4 $T=8830 1770 0 0 $X=8750 $Y=1520
X13 4 M2_M1_CDNS_5 $T=420 2020 0 90 $X=290 $Y=1940
X14 4 M2_M1_CDNS_5 $T=1680 -1770 0 90 $X=1550 $Y=-1850
X15 5 M2_M1_CDNS_5 $T=3210 -1470 0 0 $X=3130 $Y=-1600
X16 6 M2_M1_CDNS_5 $T=4220 -2030 0 180 $X=4140 $Y=-2160
X17 5 M2_M1_CDNS_5 $T=4910 -1460 0 0 $X=4830 $Y=-1590
X18 7 M2_M1_CDNS_5 $T=5310 1440 0 0 $X=5230 $Y=1310
X19 8 M2_M1_CDNS_5 $T=6360 1470 0 90 $X=6230 $Y=1390
X20 7 M2_M1_CDNS_5 $T=6800 -2140 0 90 $X=6670 $Y=-2220
X21 8 M2_M1_CDNS_5 $T=8400 1470 0 90 $X=8270 $Y=1390
X22 6 M2_M1_CDNS_5 $T=8760 -2150 0 180 $X=8680 $Y=-2280
X23 9 10 cellTmpl_CDNS_7 $T=120 -100 1 0 $X=0 $Y=-3760
X24 4 9 10 1 INV_1X_small_layout $T=0 0 0 0 $X=0 $Y=0
X25 6 9 10 5 INV_1X_small_layout $T=3800 40 1 0 $X=3800 $Y=-3760
X26 3 9 10 7 INV_1X_small_layout $T=3800 0 0 0 $X=3800 $Y=0
X27 7 9 10 8 INV_1X_small_layout $T=5200 0 0 0 $X=5200 $Y=0
X28 2 9 10 6 INV_1X_small_layout $T=7600 40 1 0 $X=7600 $Y=-3760
X29 4 9 10 5 2 12 ph1p3_clk_part $T=1400 40 1 0 $X=1400 $Y=-3760
X30 4 9 10 11 3 13 ph1p3_clk_part $T=1400 0 0 0 $X=1400 $Y=0
X31 1 9 10 7 2 14 ph1p3_clk_part $T=5200 40 1 0 $X=5200 $Y=-3760
X32 1 9 10 8 3 15 ph1p3_clk_part $T=6600 0 0 0 $X=6600 $Y=0
M0 1 4 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=780 $Y=2430 $dt=1
M1 12 4 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=2110 $Y=-2900 $dt=1
M2 13 4 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=2110 $Y=2460 $dt=1
M3 2 4 5 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=3290 $Y=-2660 $dt=1
M4 3 4 11 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=3290 $Y=2460 $dt=1
M5 5 6 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=4580 $Y=-2870 $dt=1
M6 7 3 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=4580 $Y=2430 $dt=1
M7 14 1 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=5910 $Y=-2900 $dt=1
M8 8 7 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=5980 $Y=2430 $dt=1
M9 2 1 7 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=7090 $Y=-2660 $dt=1
M10 15 1 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=7310 $Y=2460 $dt=1
M11 6 2 9 9 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=8380 $Y=-2870 $dt=1
M12 3 1 8 9 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=8490 $Y=2460 $dt=1
.ends ph1p3_DFF
