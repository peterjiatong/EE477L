* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : INV_1X_small_layout                          *
* Netlisted  : Thu Nov  7 20:00:02 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_3 D_drain_1 S_source_0 3
** N=3 EP=3 FDC=1
M0 D_drain_1 3 S_source_0 S_source_0 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_4                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_4 D_drain_1 S_source_0 3 B
** N=5 EP=4 FDC=1
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=20.6614 scb=0.0218476 scc=0.000360984 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout gnd! in out vdd!
** N=4 EP=4 FDC=2
X0 out gnd! in nmos1v_CDNS_3 $T=780 900 0 0 $X=360 $Y=700
X1 out vdd! in vdd! pmos1v_CDNS_4 $T=780 2430 0 0 $X=360 $Y=2230
.ends INV_1X_small_layout
