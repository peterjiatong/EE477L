* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph2p1_MAC                                    *
* Netlisted  : Sat Nov 23 21:11:52 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_8                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_8 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_9                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_9 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_10                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_10 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_11                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_11 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_12                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_12 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_13                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_13 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_14                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_14 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_15                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_15 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_16                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_16 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_17                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_17 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_18                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_18 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_new                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_new 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 3 M1_PO_CDNS_14 $T=1020 1750 0 90 $X=900 $Y=1650
X1 1 2 cellTmpl_CDNS_18 $T=50 150 0 0 $X=-70 $Y=10
M0 4 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.3086 scb=0.00950139 scc=0.000267597 $X=1140 $Y=930 $dt=0
.ends INV_1X_new

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_19                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_19 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_20                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_20 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_20

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_21                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_21 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_21

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X_small                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_14 $T=690 1680 0 90 $X=570 $Y=1580
X1 4 M1_PO_CDNS_14 $T=1930 1650 0 90 $X=1810 $Y=1550
X2 3 1 6 3 nmos1v_CDNS_19 $T=810 1000 0 0 $X=390 $Y=800
X3 6 4 5 3 nmos1v_CDNS_19 $T=2050 1000 0 0 $X=1630 $Y=800
X4 2 1 5 3 2 pmos1v_CDNS_20 $T=810 2440 0 0 $X=390 $Y=2240
X5 2 4 5 3 2 pmos1v_CDNS_20 $T=2050 2450 0 0 $X=1630 $Y=2250
X6 2 3 cellTmpl_CDNS_21 $T=240 210 0 0 $X=120 $Y=70
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=810 $Y=1000 $dt=0
M1 5 4 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=2050 $Y=1000 $dt=0
.ends NAND2_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6
*.DEVICECLIMB
** N=7 EP=6 FDC=3
X0 2 3 6 5 INV_1X_new $T=2480 -10 0 0 $X=2410 $Y=0
X1 1 2 3 4 6 7 NAND2_1X_small $T=-110 -70 0 0 $X=10 $Y=0
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_22                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_22 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_23                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_23 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_23

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_24                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_24 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_24

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_25                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_25 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_25

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_26                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_26 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_26

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_27                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_27 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_27

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_28                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_28 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_28

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_29                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_29 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_29

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR_small                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR_small 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=9
X0 1 M2_M1_CDNS_1 $T=350 1340 0 90 $X=220 $Y=1260
X1 6 M2_M1_CDNS_1 $T=5510 3180 0 90 $X=5380 $Y=3100
X2 6 M2_M1_CDNS_1 $T=6740 3180 0 90 $X=6610 $Y=3100
X3 1 M1_PO_CDNS_14 $T=580 1660 0 90 $X=460 $Y=1560
X4 4 M1_PO_CDNS_14 $T=1990 1480 0 90 $X=1870 $Y=1380
X5 4 M1_PO_CDNS_22 $T=5990 1680 0 90 $X=5790 $Y=1580
X6 1 M1_PO_CDNS_22 $T=7100 1350 0 90 $X=6900 $Y=1250
X7 7 M1_PO_CDNS_23 $T=3070 1660 0 90 $X=2870 $Y=1560
X8 8 M1_PO_CDNS_23 $T=4410 1540 0 90 $X=4210 $Y=1440
X9 8 M3_M2_CDNS_24 $T=1210 1540 0 90 $X=1010 $Y=1440
X10 8 M3_M2_CDNS_24 $T=4410 1540 0 90 $X=4210 $Y=1440
X11 8 M2_M1_CDNS_25 $T=1210 1540 0 90 $X=1010 $Y=1440
X12 4 M2_M1_CDNS_25 $T=1820 1880 0 90 $X=1620 $Y=1780
X13 8 M2_M1_CDNS_25 $T=4410 1540 0 90 $X=4210 $Y=1440
X14 4 M2_M1_CDNS_26 $T=5990 1680 0 90 $X=5790 $Y=1580
X15 1 M2_M1_CDNS_26 $T=7100 1350 0 90 $X=6900 $Y=1250
X16 2 3 cellTmpl_CDNS_27 $T=120 140 0 0 $X=0 $Y=0
X17 2 1 8 3 2 pmos1v_CDNS_28 $T=700 2180 0 0 $X=280 $Y=1980
X18 2 4 7 3 2 pmos1v_CDNS_28 $T=2110 2170 0 0 $X=1690 $Y=1970
X19 2 7 6 3 2 pmos1v_CDNS_28 $T=3270 2160 0 0 $X=2850 $Y=1960
X20 2 8 6 3 2 pmos1v_CDNS_28 $T=4610 2160 0 0 $X=4190 $Y=1960
X21 6 4 5 3 2 pmos1v_CDNS_28 $T=6140 2120 0 0 $X=5720 $Y=1920
X22 6 1 5 3 2 pmos1v_CDNS_28 $T=7250 2160 0 0 $X=6830 $Y=1960
X23 3 1 8 3 nmos1v_CDNS_29 $T=700 590 0 0 $X=280 $Y=390
X24 3 4 7 3 nmos1v_CDNS_29 $T=2110 580 0 0 $X=1690 $Y=380
X25 3 7 9 3 nmos1v_CDNS_29 $T=3270 580 0 0 $X=2850 $Y=380
X26 9 8 5 3 nmos1v_CDNS_29 $T=4610 580 0 0 $X=4190 $Y=380
X27 3 4 10 3 nmos1v_CDNS_29 $T=6140 600 0 0 $X=5720 $Y=400
X28 10 1 5 3 nmos1v_CDNS_29 $T=7250 650 0 0 $X=6830 $Y=450
M0 8 1 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.45462 scb=0.00478425 scc=6.8709e-05 $X=700 $Y=590 $dt=0
M1 7 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=2110 $Y=580 $dt=0
M2 9 7 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=3270 $Y=580 $dt=0
M3 5 8 9 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=4610 $Y=580 $dt=0
M4 10 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 $X=6140 $Y=600 $dt=0
M5 5 1 10 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=7250 $Y=650 $dt=0
M6 7 4 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.1869 scb=0.0086398 scc=0.00051649 $X=2110 $Y=2170 $dt=1
M7 6 7 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3270 $Y=2160 $dt=1
M8 6 8 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4610 $Y=2160 $dt=1
.ends XOR_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 8 9 13
*.DEVICECLIMB
** N=13 EP=9 FDC=12
X0 4 M3_M2_CDNS_8 $T=6750 2480 0 0 $X=6670 $Y=2230
X1 4 M3_M2_CDNS_8 $T=9120 2880 0 0 $X=9040 $Y=2630
X2 4 M2_M1_CDNS_16 $T=6750 2480 0 0 $X=6670 $Y=2230
X3 4 M2_M1_CDNS_16 $T=9120 2880 0 0 $X=9040 $Y=2630
X4 4 M1_PO_CDNS_17 $T=6750 2480 0 0 $X=6650 $Y=2230
X5 4 M1_PO_CDNS_17 $T=9120 2880 0 0 $X=9020 $Y=2630
X6 1 3 2 4 6 9 AND $T=7790 0 0 0 $X=7800 $Y=0
X7 1 3 2 4 5 13 7 8 10 11 XOR_small $T=0 0 0 0 $X=0 $Y=0
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_33                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_33 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_33

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_1X_small                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=-310 120 0 0 $X=-430 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1000 $Y=830 $dt=0
M1 4 5 6 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1210 $Y=830 $dt=0
.ends NAND_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_2X_small1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_2X_small1 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=130 160 0 0 $X=10 $Y=20
M0 6 4 2 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=7.66878 scb=0.00580736 scc=7.77234e-05 $X=940 $Y=890 $dt=0
M1 3 5 6 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=11.676 scb=0.0124835 scc=0.000479408 $X=940 $Y=1100 $dt=0
.ends NAND_2X_small1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_39                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_39 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_39

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR1 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=6
X0 6 M2_M1_CDNS_1 $T=1210 1480 0 90 $X=1080 $Y=1400
X1 7 M2_M1_CDNS_1 $T=2250 1860 0 90 $X=2120 $Y=1780
X2 6 M2_M1_CDNS_1 $T=2950 1480 0 90 $X=2820 $Y=1400
X3 8 M2_M1_CDNS_1 $T=3370 650 0 0 $X=3290 $Y=520
X4 9 M2_M1_CDNS_1 $T=3370 3080 0 0 $X=3290 $Y=2950
X5 9 M2_M1_CDNS_1 $T=3930 3080 0 0 $X=3850 $Y=2950
X6 7 M2_M1_CDNS_1 $T=4680 1860 0 90 $X=4550 $Y=1780
X7 9 M2_M1_CDNS_1 $T=4890 3070 0 0 $X=4810 $Y=2940
X8 8 M2_M1_CDNS_1 $T=5840 640 0 0 $X=5760 $Y=510
X9 9 M2_M1_CDNS_1 $T=6260 3080 0 0 $X=6180 $Y=2950
X10 6 M1_PO_CDNS_14 $T=4020 1500 0 90 $X=3900 $Y=1400
X11 7 M1_PO_CDNS_14 $T=5020 1730 0 90 $X=4900 $Y=1630
X12 2 3 6 2 nmos1v_CDNS_19 $T=830 840 0 0 $X=410 $Y=640
X13 2 4 7 2 nmos1v_CDNS_19 $T=1790 840 0 0 $X=1370 $Y=640
X14 1 3 6 2 1 pmos1v_CDNS_20 $T=830 2320 0 0 $X=410 $Y=2120
X15 1 4 7 2 1 pmos1v_CDNS_20 $T=1790 2320 0 0 $X=1370 $Y=2120
X16 1 4 9 2 1 pmos1v_CDNS_28 $T=3120 2080 0 0 $X=2700 $Y=1880
X17 9 6 5 2 1 pmos1v_CDNS_28 $T=4090 2140 0 0 $X=3670 $Y=1940
X18 9 7 5 2 1 pmos1v_CDNS_28 $T=5050 2140 0 0 $X=4630 $Y=1940
X19 1 3 9 2 1 pmos1v_CDNS_28 $T=6010 2140 0 0 $X=5590 $Y=1940
X20 2 4 8 2 nmos1v_CDNS_29 $T=3120 780 0 0 $X=2700 $Y=580
X21 10 6 5 2 nmos1v_CDNS_29 $T=4090 760 0 0 $X=3670 $Y=560
X22 10 7 2 2 nmos1v_CDNS_29 $T=5050 770 0 0 $X=4630 $Y=570
X23 8 3 5 2 nmos1v_CDNS_29 $T=6010 770 0 0 $X=5590 $Y=570
X24 1 2 cellTmpl_CDNS_39 $T=180 120 0 0 $X=60 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=830 $Y=840 $dt=0
M1 7 4 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1790 $Y=840 $dt=0
M2 8 4 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=3120 $Y=780 $dt=0
M3 5 6 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4126 scb=0.0095497 scc=0.000351079 $X=4090 $Y=760 $dt=0
M4 2 7 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=5050 $Y=770 $dt=0
M5 5 3 8 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=6010 $Y=770 $dt=0
.ends XOR1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder1_small                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder1_small 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 22 23
*.DEVICECLIMB
** N=23 EP=16 FDC=18
X0 8 M2_M1_CDNS_1 $T=6580 1900 0 0 $X=6500 $Y=1770
X1 9 M2_M1_CDNS_1 $T=15190 1730 0 90 $X=15060 $Y=1650
X2 8 M3_M2_CDNS_2 $T=6970 950 0 0 $X=6890 $Y=820
X3 8 M3_M2_CDNS_2 $T=14100 570 0 90 $X=13970 $Y=490
X4 1 M3_M2_CDNS_8 $T=590 2080 0 90 $X=340 $Y=2000
X5 3 M3_M2_CDNS_8 $T=2300 3150 0 90 $X=2050 $Y=3070
X6 1 M3_M2_CDNS_8 $T=17380 1890 0 0 $X=17300 $Y=1640
X7 3 M3_M2_CDNS_8 $T=19040 3010 0 0 $X=18960 $Y=2760
X8 8 M1_PO_CDNS_13 $T=8510 1970 0 0 $X=8410 $Y=1720
X9 8 M1_PO_CDNS_13 $T=16110 1570 0 0 $X=16010 $Y=1320
X10 9 M1_PO_CDNS_13 $T=20260 1840 0 0 $X=20160 $Y=1590
X11 1 M1_PO_CDNS_14 $T=690 1610 0 0 $X=590 $Y=1490
X12 3 M1_PO_CDNS_14 $T=1650 1990 0 0 $X=1550 $Y=1870
X13 5 M1_PO_CDNS_14 $T=7590 1960 0 0 $X=7490 $Y=1840
X14 10 M1_PO_CDNS_14 $T=19320 1680 0 0 $X=19220 $Y=1560
X15 8 M2_M1_CDNS_15 $T=8510 1970 0 0 $X=8430 $Y=1720
X16 8 M2_M1_CDNS_15 $T=16110 1570 0 0 $X=16030 $Y=1320
X17 9 M2_M1_CDNS_15 $T=20260 1840 0 0 $X=20180 $Y=1590
X18 1 M2_M1_CDNS_16 $T=590 2080 0 90 $X=340 $Y=2000
X19 3 M2_M1_CDNS_16 $T=2300 3150 0 90 $X=2050 $Y=3070
X20 1 M2_M1_CDNS_16 $T=17380 1890 0 0 $X=17300 $Y=1640
X21 3 M2_M1_CDNS_16 $T=19040 3010 0 0 $X=18960 $Y=2760
X22 1 M1_PO_CDNS_17 $T=590 2080 0 90 $X=340 $Y=1980
X23 3 M1_PO_CDNS_17 $T=2300 3150 0 90 $X=2050 $Y=3050
X24 1 M1_PO_CDNS_17 $T=17380 1890 0 0 $X=17280 $Y=1640
X25 3 M1_PO_CDNS_17 $T=19040 3010 0 0 $X=18940 $Y=2760
X26 2 4 1 10 3 20 NAND_1X_small $T=16970 30 0 0 $X=16540 $Y=10
X27 2 4 9 7 10 21 NAND_1X_small $T=19810 30 0 0 $X=19380 $Y=10
X28 2 4 9 5 8 19 NAND_2X_small1 $T=13690 -10 0 0 $X=13700 $Y=10
X29 2 4 1 3 8 11 12 15 22 16 XOR1 $T=-40 30 0 0 $X=20 $Y=10
X30 2 4 5 8 6 13 14 17 23 18 XOR1 $T=6800 30 0 0 $X=6860 $Y=10
.ends full_adder1_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: multiplier                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt multiplier 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
** N=238 EP=50 FDC=456
X0 2 M2_M1_CDNS_1 $T=170 4730 0 0 $X=90 $Y=4600
X1 2 M2_M1_CDNS_1 $T=180 890 0 0 $X=100 $Y=760
X2 19 M2_M1_CDNS_1 $T=4340 11800 0 0 $X=4260 $Y=11670
X3 20 M2_M1_CDNS_1 $T=8880 12210 0 0 $X=8800 $Y=12080
X4 21 M2_M1_CDNS_1 $T=13420 4530 0 0 $X=13340 $Y=4400
X5 22 M2_M1_CDNS_1 $T=17560 15460 0 0 $X=17480 $Y=15330
X6 23 M2_M1_CDNS_1 $T=21930 4780 0 0 $X=21850 $Y=4650
X7 24 M2_M1_CDNS_1 $T=29730 11900 0 0 $X=29650 $Y=11770
X8 25 M2_M1_CDNS_1 $T=31310 15530 0 0 $X=31230 $Y=15400
X9 26 M2_M1_CDNS_1 $T=35410 9580 0 0 $X=35330 $Y=9450
X10 27 M2_M1_CDNS_1 $T=41980 11840 0 0 $X=41900 $Y=11710
X11 28 M2_M1_CDNS_1 $T=43890 4790 0 0 $X=43810 $Y=4660
X12 29 M3_M2_CDNS_2 $T=4340 13390 0 0 $X=4260 $Y=13260
X13 30 M3_M2_CDNS_2 $T=7370 12440 0 0 $X=7290 $Y=12310
X14 30 M3_M2_CDNS_2 $T=8600 9080 0 0 $X=8520 $Y=8950
X15 8 M3_M2_CDNS_2 $T=10370 18740 0 0 $X=10290 $Y=18610
X16 31 M3_M2_CDNS_2 $T=13190 12020 0 0 $X=13110 $Y=11890
X17 23 M3_M2_CDNS_2 $T=19690 2880 0 90 $X=19560 $Y=2800
X18 32 M3_M2_CDNS_2 $T=26840 17540 0 90 $X=26710 $Y=17460
X19 33 M3_M2_CDNS_2 $T=35760 21100 0 0 $X=35680 $Y=20970
X20 1 M4_M3_CDNS_3 $T=1390 19500 0 0 $X=1310 $Y=19250
X21 29 M4_M3_CDNS_3 $T=3370 8280 0 0 $X=3290 $Y=8030
X22 7 M4_M3_CDNS_3 $T=4510 16920 0 0 $X=4430 $Y=16670
X23 19 M4_M3_CDNS_3 $T=5400 9800 0 0 $X=5320 $Y=9550
X24 7 M4_M3_CDNS_3 $T=7950 19550 0 0 $X=7870 $Y=19300
X25 34 M4_M3_CDNS_3 $T=8750 8160 0 0 $X=8670 $Y=7910
X26 35 M4_M3_CDNS_3 $T=10750 19470 0 0 $X=10670 $Y=19220
X27 36 M4_M3_CDNS_3 $T=11680 11800 0 0 $X=11600 $Y=11550
X28 31 M4_M3_CDNS_3 $T=12950 9830 0 0 $X=12870 $Y=9580
X29 11 M4_M3_CDNS_3 $T=13290 16990 0 0 $X=13210 $Y=16740
X30 21 M4_M3_CDNS_3 $T=14070 2580 0 90 $X=13820 $Y=2500
X31 20 M4_M3_CDNS_3 $T=15700 9710 0 0 $X=15620 $Y=9460
X32 36 M4_M3_CDNS_3 $T=22150 6400 0 0 $X=22070 $Y=6150
X33 20 M4_M3_CDNS_3 $T=24490 750 0 0 $X=24410 $Y=500
X34 11 M4_M3_CDNS_3 $T=25590 19380 0 0 $X=25510 $Y=19130
X35 32 M4_M3_CDNS_3 $T=25970 20660 0 0 $X=25890 $Y=20410
X36 37 M4_M3_CDNS_3 $T=26370 19410 0 0 $X=26290 $Y=19160
X37 38 M4_M3_CDNS_3 $T=26600 23000 0 0 $X=26520 $Y=22750
X38 24 M4_M3_CDNS_3 $T=28540 8430 0 0 $X=28460 $Y=8180
X39 24 M4_M3_CDNS_3 $T=28700 9810 0 0 $X=28620 $Y=9560
X40 39 M4_M3_CDNS_3 $T=29280 19170 0 0 $X=29200 $Y=18920
X41 28 M4_M3_CDNS_3 $T=35970 2380 0 0 $X=35890 $Y=2130
X42 40 M4_M3_CDNS_3 $T=38260 18710 0 0 $X=38180 $Y=18460
X43 39 M4_M3_CDNS_3 $T=39640 17490 0 0 $X=39560 $Y=17240
X44 28 M4_M3_CDNS_3 $T=42090 2930 0 90 $X=41840 $Y=2850
X45 41 M4_M3_CDNS_3 $T=43850 8260 0 0 $X=43770 $Y=8010
X46 42 M4_M3_CDNS_3 $T=43880 660 0 0 $X=43800 $Y=410
X47 40 M4_M3_CDNS_3 $T=46340 18970 0 0 $X=46260 $Y=18720
X48 38 M4_M3_CDNS_4 $T=34850 16990 0 0 $X=34770 $Y=16740
X49 1 M4_M3_CDNS_5 $T=1390 21140 0 0 $X=1310 $Y=21010
X50 29 M4_M3_CDNS_5 $T=3650 6110 0 0 $X=3570 $Y=5980
X51 19 M4_M3_CDNS_5 $T=6680 2460 0 0 $X=6600 $Y=2330
X52 32 M4_M3_CDNS_5 $T=13170 22790 0 0 $X=13090 $Y=22660
X53 31 M4_M3_CDNS_5 $T=13680 4950 0 0 $X=13600 $Y=4820
X54 11 M4_M3_CDNS_5 $T=14530 13310 0 0 $X=14450 $Y=13180
X55 11 M4_M3_CDNS_5 $T=14530 15600 0 0 $X=14450 $Y=15470
X56 21 M4_M3_CDNS_5 $T=21870 1570 0 0 $X=21790 $Y=1440
X57 34 M4_M3_CDNS_5 $T=23120 3950 0 0 $X=23040 $Y=3820
X58 37 M4_M3_CDNS_5 $T=28320 12210 0 0 $X=28240 $Y=12080
X59 42 M4_M3_CDNS_5 $T=28540 230 0 90 $X=28410 $Y=150
X60 41 M4_M3_CDNS_5 $T=28550 7610 0 90 $X=28420 $Y=7530
X61 35 M4_M3_CDNS_5 $T=33860 19960 0 90 $X=33730 $Y=19880
X62 1 M3_M2_CDNS_6 $T=1390 21140 0 0 $X=1310 $Y=20890
X63 7 M3_M2_CDNS_6 $T=4510 16920 0 0 $X=4430 $Y=16670
X64 34 M3_M2_CDNS_6 $T=8750 8160 0 0 $X=8670 $Y=7910
X65 35 M3_M2_CDNS_6 $T=10750 19470 0 0 $X=10670 $Y=19220
X66 36 M3_M2_CDNS_6 $T=11680 11800 0 0 $X=11600 $Y=11550
X67 32 M3_M2_CDNS_6 $T=13170 22790 0 0 $X=13090 $Y=22540
X68 11 M3_M2_CDNS_6 $T=13290 16990 0 0 $X=13210 $Y=16740
X69 11 M3_M2_CDNS_6 $T=14530 13310 0 0 $X=14450 $Y=13060
X70 11 M3_M2_CDNS_6 $T=14530 15600 0 0 $X=14450 $Y=15350
X71 36 M3_M2_CDNS_6 $T=22150 6400 0 0 $X=22070 $Y=6150
X72 20 M3_M2_CDNS_6 $T=24490 750 0 0 $X=24410 $Y=500
X73 37 M3_M2_CDNS_6 $T=26370 19410 0 0 $X=26290 $Y=19160
X74 38 M3_M2_CDNS_6 $T=26600 23000 0 0 $X=26520 $Y=22750
X75 43 M3_M2_CDNS_6 $T=28820 19250 0 0 $X=28740 $Y=19000
X76 39 M3_M2_CDNS_6 $T=29280 19170 0 0 $X=29200 $Y=18920
X77 35 M3_M2_CDNS_6 $T=33860 19960 0 90 $X=33610 $Y=19880
X78 43 M3_M2_CDNS_6 $T=34220 19150 0 0 $X=34140 $Y=18900
X79 28 M3_M2_CDNS_6 $T=35970 2380 0 0 $X=35890 $Y=2130
X80 39 M3_M2_CDNS_6 $T=39640 17490 0 0 $X=39560 $Y=17240
X81 41 M3_M2_CDNS_6 $T=43850 8260 0 0 $X=43770 $Y=8010
X82 42 M3_M2_CDNS_6 $T=43880 660 0 0 $X=43800 $Y=410
X83 40 M3_M2_CDNS_6 $T=46340 18970 0 0 $X=46260 $Y=18720
X84 1 M3_M2_CDNS_7 $T=1390 19500 0 0 $X=1310 $Y=19250
X85 29 M3_M2_CDNS_7 $T=3370 8280 0 0 $X=3290 $Y=8030
X86 19 M3_M2_CDNS_7 $T=5400 9800 0 0 $X=5320 $Y=9550
X87 7 M3_M2_CDNS_7 $T=7950 19550 0 0 $X=7870 $Y=19300
X88 31 M3_M2_CDNS_7 $T=12950 9830 0 0 $X=12870 $Y=9580
X89 21 M3_M2_CDNS_7 $T=14070 2580 0 90 $X=13820 $Y=2500
X90 20 M3_M2_CDNS_7 $T=15700 9710 0 0 $X=15620 $Y=9460
X91 11 M3_M2_CDNS_7 $T=25590 19380 0 0 $X=25510 $Y=19130
X92 32 M3_M2_CDNS_7 $T=25970 20660 0 0 $X=25890 $Y=20410
X93 24 M3_M2_CDNS_7 $T=28540 8430 0 0 $X=28460 $Y=8180
X94 24 M3_M2_CDNS_7 $T=28700 9810 0 0 $X=28620 $Y=9560
X95 40 M3_M2_CDNS_7 $T=38260 18710 0 0 $X=38180 $Y=18460
X96 28 M3_M2_CDNS_7 $T=42090 2930 0 90 $X=41840 $Y=2850
X97 2 M3_M2_CDNS_8 $T=160 15480 0 0 $X=80 $Y=15230
X98 2 M3_M2_CDNS_8 $T=160 21130 0 0 $X=80 $Y=20880
X99 2 M3_M2_CDNS_8 $T=170 9270 0 0 $X=90 $Y=9020
X100 2 M3_M2_CDNS_8 $T=170 13790 0 0 $X=90 $Y=13540
X101 44 M3_M2_CDNS_8 $T=500 8210 0 0 $X=420 $Y=7960
X102 1 M3_M2_CDNS_8 $T=1350 15570 0 0 $X=1270 $Y=15320
X103 1 M3_M2_CDNS_8 $T=1360 13320 0 0 $X=1280 $Y=13070
X104 45 M3_M2_CDNS_8 $T=4380 23070 0 90 $X=4130 $Y=22990
X105 29 M3_M2_CDNS_8 $T=4340 15320 0 0 $X=4260 $Y=15070
X106 30 M3_M2_CDNS_8 $T=5400 21130 0 0 $X=5320 $Y=20880
X107 7 M3_M2_CDNS_8 $T=5740 15570 0 0 $X=5660 $Y=15320
X108 7 M3_M2_CDNS_8 $T=5750 13320 0 0 $X=5670 $Y=13070
X109 44 M3_M2_CDNS_8 $T=6590 5910 0 0 $X=6510 $Y=5660
X110 46 M3_M2_CDNS_8 $T=7520 22860 0 0 $X=7440 $Y=22610
X111 46 M3_M2_CDNS_8 $T=7960 21030 0 0 $X=7880 $Y=20780
X112 47 M3_M2_CDNS_8 $T=8730 15340 0 0 $X=8650 $Y=15090
X113 8 M3_M2_CDNS_8 $T=8980 17010 0 0 $X=8900 $Y=16760
X114 8 M3_M2_CDNS_8 $T=10140 15570 0 0 $X=10060 $Y=15320
X115 8 M3_M2_CDNS_8 $T=10150 13320 0 0 $X=10070 $Y=13070
X116 31 M3_M2_CDNS_8 $T=12100 19160 0 0 $X=12020 $Y=18910
X117 45 M3_M2_CDNS_8 $T=12260 20780 0 0 $X=12180 $Y=20530
X118 48 M3_M2_CDNS_8 $T=13150 15340 0 0 $X=13070 $Y=15090
X119 49 M3_M2_CDNS_8 $T=14690 20780 0 0 $X=14610 $Y=20530
X120 41 M3_M2_CDNS_8 $T=15670 8330 0 0 $X=15590 $Y=8080
X121 42 M3_M2_CDNS_8 $T=16600 750 0 0 $X=16520 $Y=500
X122 49 M3_M2_CDNS_8 $T=17570 22850 0 0 $X=17490 $Y=22600
X123 43 M3_M2_CDNS_8 $T=22230 22840 0 0 $X=22150 $Y=22590
X124 43 M3_M2_CDNS_8 $T=28820 20830 0 0 $X=28740 $Y=20580
X125 33 M3_M2_CDNS_8 $T=35370 22940 0 0 $X=35290 $Y=22690
X126 2 M2_M1_CDNS_9 $T=160 15480 0 0 $X=80 $Y=15230
X127 2 M2_M1_CDNS_9 $T=160 21130 0 0 $X=80 $Y=20880
X128 2 M2_M1_CDNS_9 $T=170 9270 0 0 $X=90 $Y=9020
X129 2 M2_M1_CDNS_9 $T=170 13790 0 0 $X=90 $Y=13540
X130 44 M2_M1_CDNS_9 $T=500 8210 0 0 $X=420 $Y=7960
X131 45 M2_M1_CDNS_9 $T=4380 23070 0 90 $X=4130 $Y=22990
X132 29 M2_M1_CDNS_9 $T=4340 15320 0 0 $X=4260 $Y=15070
X133 30 M2_M1_CDNS_9 $T=5400 21130 0 0 $X=5320 $Y=20880
X134 47 M2_M1_CDNS_9 $T=8730 15340 0 0 $X=8650 $Y=15090
X135 31 M2_M1_CDNS_9 $T=12100 19160 0 0 $X=12020 $Y=18910
X136 48 M2_M1_CDNS_9 $T=13150 15340 0 0 $X=13070 $Y=15090
X137 49 M2_M1_CDNS_9 $T=17570 22850 0 0 $X=17490 $Y=22600
X138 43 M2_M1_CDNS_9 $T=22230 22840 0 0 $X=22150 $Y=22590
X139 43 M2_M1_CDNS_9 $T=28820 20830 0 0 $X=28740 $Y=20580
X140 33 M2_M1_CDNS_9 $T=35370 22940 0 0 $X=35290 $Y=22690
X141 40 M2_M1_CDNS_9 $T=46340 18970 0 0 $X=46260 $Y=18720
X142 43 M5_M4_CDNS_10 $T=34220 19150 0 0 $X=34140 $Y=18900
X143 38 M5_M4_CDNS_10 $T=34850 16990 0 0 $X=34770 $Y=16740
X144 43 M4_M3_CDNS_11 $T=28820 19250 0 0 $X=28740 $Y=19000
X145 43 M4_M3_CDNS_11 $T=34220 19150 0 0 $X=34140 $Y=18900
X146 43 M5_M4_CDNS_12 $T=28820 19250 0 0 $X=28740 $Y=19120
X147 38 M5_M4_CDNS_12 $T=35550 19590 0 0 $X=35470 $Y=19460
X148 1 M1_PO_CDNS_13 $T=1390 17230 0 0 $X=1290 $Y=16980
X149 1 M1_PO_CDNS_13 $T=1390 24660 0 0 $X=1290 $Y=24410
X150 3 M1_PO_CDNS_13 $T=2770 22320 0 90 $X=2520 $Y=22220
X151 5 M1_PO_CDNS_13 $T=2650 13610 0 0 $X=2550 $Y=13360
X152 4 M1_PO_CDNS_13 $T=2750 17050 0 0 $X=2650 $Y=16800
X153 1 M1_PO_CDNS_13 $T=4410 23850 0 0 $X=4310 $Y=23600
X154 4 M1_PO_CDNS_13 $T=5790 16970 0 0 $X=5690 $Y=16720
X155 9 M1_PO_CDNS_13 $T=7290 23970 0 90 $X=7040 $Y=23870
X156 5 M1_PO_CDNS_13 $T=7180 13450 0 0 $X=7080 $Y=13200
X157 3 M1_PO_CDNS_13 $T=8720 22330 0 90 $X=8470 $Y=22230
X158 3 M1_PO_CDNS_13 $T=9910 24890 0 90 $X=9660 $Y=24790
X159 4 M1_PO_CDNS_13 $T=10210 17010 0 0 $X=10110 $Y=16760
X160 7 M1_PO_CDNS_13 $T=11550 22710 0 0 $X=11450 $Y=22460
X161 5 M1_PO_CDNS_13 $T=11730 13390 0 0 $X=11630 $Y=13140
X162 9 M1_PO_CDNS_13 $T=13230 23970 0 90 $X=12980 $Y=23870
X163 4 M1_PO_CDNS_13 $T=14630 17040 0 0 $X=14530 $Y=16790
X164 7 M1_PO_CDNS_13 $T=15790 22330 0 90 $X=15540 $Y=22230
X165 5 M1_PO_CDNS_13 $T=15980 13520 0 0 $X=15880 $Y=13270
X166 3 M1_PO_CDNS_13 $T=17780 24480 0 0 $X=17680 $Y=24230
X167 8 M1_PO_CDNS_13 $T=20560 22320 0 90 $X=20310 $Y=22220
X168 9 M1_PO_CDNS_13 $T=22240 23950 0 0 $X=22140 $Y=23700
X169 8 M1_PO_CDNS_13 $T=24880 22320 0 90 $X=24630 $Y=22220
X170 3 M1_PO_CDNS_13 $T=26710 24400 0 0 $X=26610 $Y=24150
X171 24 M1_PO_CDNS_13 $T=28540 6330 0 0 $X=28440 $Y=6080
X172 11 M1_PO_CDNS_13 $T=29350 22530 0 0 $X=29250 $Y=22280
X173 22 M1_PO_CDNS_13 $T=29800 13490 0 0 $X=29700 $Y=13240
X174 9 M1_PO_CDNS_13 $T=31140 23850 0 0 $X=31040 $Y=23600
X175 25 M1_PO_CDNS_13 $T=31170 13680 0 0 $X=31070 $Y=13430
X176 40 M1_PO_CDNS_13 $T=31860 16950 0 0 $X=31760 $Y=16700
X177 11 M1_PO_CDNS_13 $T=33650 22300 0 90 $X=33400 $Y=22200
X178 27 M1_PO_CDNS_13 $T=35890 9730 0 0 $X=35790 $Y=9480
X179 1 M2_M1_CDNS_15 $T=1390 17230 0 0 $X=1310 $Y=16980
X180 1 M2_M1_CDNS_15 $T=1390 24660 0 0 $X=1310 $Y=24410
X181 3 M2_M1_CDNS_15 $T=2770 22320 0 90 $X=2520 $Y=22240
X182 5 M2_M1_CDNS_15 $T=2650 13610 0 0 $X=2570 $Y=13360
X183 4 M2_M1_CDNS_15 $T=2750 17050 0 0 $X=2670 $Y=16800
X184 1 M2_M1_CDNS_15 $T=4410 23850 0 0 $X=4330 $Y=23600
X185 4 M2_M1_CDNS_15 $T=5790 16970 0 0 $X=5710 $Y=16720
X186 9 M2_M1_CDNS_15 $T=7290 23970 0 90 $X=7040 $Y=23890
X187 5 M2_M1_CDNS_15 $T=7180 13450 0 0 $X=7100 $Y=13200
X188 3 M2_M1_CDNS_15 $T=8720 22330 0 90 $X=8470 $Y=22250
X189 3 M2_M1_CDNS_15 $T=9910 24890 0 90 $X=9660 $Y=24810
X190 4 M2_M1_CDNS_15 $T=10210 17010 0 0 $X=10130 $Y=16760
X191 7 M2_M1_CDNS_15 $T=11550 22710 0 0 $X=11470 $Y=22460
X192 5 M2_M1_CDNS_15 $T=11730 13390 0 0 $X=11650 $Y=13140
X193 9 M2_M1_CDNS_15 $T=13230 23970 0 90 $X=12980 $Y=23890
X194 4 M2_M1_CDNS_15 $T=14630 17040 0 0 $X=14550 $Y=16790
X195 7 M2_M1_CDNS_15 $T=15790 22330 0 90 $X=15540 $Y=22250
X196 5 M2_M1_CDNS_15 $T=15980 13520 0 0 $X=15900 $Y=13270
X197 3 M2_M1_CDNS_15 $T=17780 24480 0 0 $X=17700 $Y=24230
X198 8 M2_M1_CDNS_15 $T=20560 22320 0 90 $X=20310 $Y=22240
X199 9 M2_M1_CDNS_15 $T=22240 23950 0 0 $X=22160 $Y=23700
X200 8 M2_M1_CDNS_15 $T=24880 22320 0 90 $X=24630 $Y=22240
X201 3 M2_M1_CDNS_15 $T=26710 24400 0 0 $X=26630 $Y=24150
X202 24 M2_M1_CDNS_15 $T=28540 6330 0 0 $X=28460 $Y=6080
X203 11 M2_M1_CDNS_15 $T=29350 22530 0 0 $X=29270 $Y=22280
X204 22 M2_M1_CDNS_15 $T=29800 13490 0 0 $X=29720 $Y=13240
X205 9 M2_M1_CDNS_15 $T=31140 23850 0 0 $X=31060 $Y=23600
X206 25 M2_M1_CDNS_15 $T=31170 13680 0 0 $X=31090 $Y=13430
X207 40 M2_M1_CDNS_15 $T=31860 16950 0 0 $X=31780 $Y=16700
X208 11 M2_M1_CDNS_15 $T=33650 22300 0 90 $X=33400 $Y=22220
X209 27 M2_M1_CDNS_15 $T=35890 9730 0 0 $X=35810 $Y=9480
X210 1 M2_M1_CDNS_16 $T=1350 15570 0 0 $X=1270 $Y=15320
X211 1 M2_M1_CDNS_16 $T=1360 13320 0 0 $X=1280 $Y=13070
X212 1 M2_M1_CDNS_16 $T=1390 21140 0 0 $X=1310 $Y=20890
X213 7 M2_M1_CDNS_16 $T=4510 16920 0 0 $X=4430 $Y=16670
X214 7 M2_M1_CDNS_16 $T=5740 15570 0 0 $X=5660 $Y=15320
X215 7 M2_M1_CDNS_16 $T=5750 13320 0 0 $X=5670 $Y=13070
X216 44 M2_M1_CDNS_16 $T=6590 5910 0 0 $X=6510 $Y=5660
X217 46 M2_M1_CDNS_16 $T=7520 22860 0 0 $X=7440 $Y=22610
X218 46 M2_M1_CDNS_16 $T=7960 21030 0 0 $X=7880 $Y=20780
X219 34 M2_M1_CDNS_16 $T=8750 8160 0 0 $X=8670 $Y=7910
X220 8 M2_M1_CDNS_16 $T=8980 17010 0 0 $X=8900 $Y=16760
X221 8 M2_M1_CDNS_16 $T=10140 15570 0 0 $X=10060 $Y=15320
X222 8 M2_M1_CDNS_16 $T=10150 13320 0 0 $X=10070 $Y=13070
X223 8 M2_M1_CDNS_16 $T=10370 18740 0 0 $X=10290 $Y=18490
X224 35 M2_M1_CDNS_16 $T=10750 19470 0 0 $X=10670 $Y=19220
X225 36 M2_M1_CDNS_16 $T=11680 11800 0 0 $X=11600 $Y=11550
X226 45 M2_M1_CDNS_16 $T=12260 20780 0 0 $X=12180 $Y=20530
X227 32 M2_M1_CDNS_16 $T=13170 22790 0 0 $X=13090 $Y=22540
X228 11 M2_M1_CDNS_16 $T=13290 16990 0 0 $X=13210 $Y=16740
X229 11 M2_M1_CDNS_16 $T=14530 13310 0 0 $X=14450 $Y=13060
X230 11 M2_M1_CDNS_16 $T=14530 15600 0 0 $X=14450 $Y=15350
X231 49 M2_M1_CDNS_16 $T=14690 20780 0 0 $X=14610 $Y=20530
X232 41 M2_M1_CDNS_16 $T=15670 8330 0 0 $X=15590 $Y=8080
X233 42 M2_M1_CDNS_16 $T=16600 750 0 0 $X=16520 $Y=500
X234 36 M2_M1_CDNS_16 $T=22150 6400 0 0 $X=22070 $Y=6150
X235 20 M2_M1_CDNS_16 $T=24490 750 0 0 $X=24410 $Y=500
X236 37 M2_M1_CDNS_16 $T=26370 19410 0 0 $X=26290 $Y=19160
X237 38 M2_M1_CDNS_16 $T=26600 23000 0 0 $X=26520 $Y=22750
X238 43 M2_M1_CDNS_16 $T=28820 19250 0 0 $X=28740 $Y=19000
X239 39 M2_M1_CDNS_16 $T=29280 19170 0 0 $X=29200 $Y=18920
X240 35 M2_M1_CDNS_16 $T=33860 19960 0 90 $X=33610 $Y=19880
X241 43 M2_M1_CDNS_16 $T=34220 19150 0 0 $X=34140 $Y=18900
X242 33 M2_M1_CDNS_16 $T=35760 21100 0 0 $X=35680 $Y=20850
X243 28 M2_M1_CDNS_16 $T=35970 2380 0 0 $X=35890 $Y=2130
X244 39 M2_M1_CDNS_16 $T=39640 17490 0 0 $X=39560 $Y=17240
X245 41 M2_M1_CDNS_16 $T=43850 8260 0 0 $X=43770 $Y=8010
X246 42 M2_M1_CDNS_16 $T=43880 660 0 0 $X=43800 $Y=410
X247 1 M1_PO_CDNS_17 $T=1350 15570 0 0 $X=1250 $Y=15320
X248 1 M1_PO_CDNS_17 $T=1360 13320 0 0 $X=1260 $Y=13070
X249 7 M1_PO_CDNS_17 $T=4510 16920 0 0 $X=4410 $Y=16670
X250 7 M1_PO_CDNS_17 $T=5740 15570 0 0 $X=5640 $Y=15320
X251 7 M1_PO_CDNS_17 $T=5750 13320 0 0 $X=5650 $Y=13070
X252 44 M1_PO_CDNS_17 $T=6590 5910 0 0 $X=6490 $Y=5660
X253 46 M1_PO_CDNS_17 $T=7520 22860 0 0 $X=7420 $Y=22610
X254 46 M1_PO_CDNS_17 $T=7960 21030 0 0 $X=7860 $Y=20780
X255 8 M1_PO_CDNS_17 $T=8980 17010 0 0 $X=8880 $Y=16760
X256 8 M1_PO_CDNS_17 $T=10140 15570 0 0 $X=10040 $Y=15320
X257 8 M1_PO_CDNS_17 $T=10150 13320 0 0 $X=10050 $Y=13070
X258 8 M1_PO_CDNS_17 $T=10370 18740 0 0 $X=10270 $Y=18490
X259 35 M1_PO_CDNS_17 $T=10750 19470 0 0 $X=10650 $Y=19220
X260 45 M1_PO_CDNS_17 $T=12260 20780 0 0 $X=12160 $Y=20530
X261 11 M1_PO_CDNS_17 $T=13290 16990 0 0 $X=13190 $Y=16740
X262 11 M1_PO_CDNS_17 $T=14530 13310 0 0 $X=14430 $Y=13060
X263 11 M1_PO_CDNS_17 $T=14530 15600 0 0 $X=14430 $Y=15350
X264 49 M1_PO_CDNS_17 $T=14690 20780 0 0 $X=14590 $Y=20530
X265 41 M1_PO_CDNS_17 $T=15670 8330 0 0 $X=15570 $Y=8080
X266 42 M1_PO_CDNS_17 $T=16600 750 0 0 $X=16500 $Y=500
X267 36 M1_PO_CDNS_17 $T=22150 6400 0 0 $X=22050 $Y=6150
X268 20 M1_PO_CDNS_17 $T=24490 750 0 0 $X=24390 $Y=500
X269 39 M1_PO_CDNS_17 $T=29280 19170 0 0 $X=29180 $Y=18920
X270 43 M1_PO_CDNS_17 $T=34220 19150 0 0 $X=34120 $Y=18900
X271 33 M1_PO_CDNS_17 $T=35760 21100 0 0 $X=35660 $Y=20850
X272 28 M1_PO_CDNS_17 $T=35970 2380 0 0 $X=35870 $Y=2130
X273 1 6 2 5 19 77 AND $T=40 14460 1 0 $X=50 $Y=10660
X274 1 6 2 4 29 76 AND $T=40 14420 0 0 $X=50 $Y=14420
X275 1 6 2 3 45 75 AND $T=40 21740 0 0 $X=50 $Y=21740
X276 7 6 2 5 20 80 AND $T=4440 14460 1 0 $X=4450 $Y=10660
X277 7 6 2 4 47 79 AND $T=4440 14420 0 0 $X=4450 $Y=14420
X278 1 6 2 9 46 78 AND $T=4440 21740 0 0 $X=4450 $Y=21740
X279 8 6 2 5 36 83 AND $T=8840 14460 1 0 $X=8850 $Y=10660
X280 8 6 2 4 48 82 AND $T=8840 14420 0 0 $X=8850 $Y=14420
X281 3 6 2 7 32 81 AND $T=8840 21740 0 0 $X=8850 $Y=21740
X282 11 6 2 5 50 93 AND $T=13240 14460 1 0 $X=13250 $Y=10660
X283 11 6 2 4 22 92 AND $T=13240 14420 0 0 $X=13250 $Y=14420
X284 9 6 2 7 49 91 AND $T=13240 21740 0 0 $X=13250 $Y=21740
X285 3 6 2 8 43 104 AND $T=17880 21740 0 0 $X=17890 $Y=21740
X286 9 6 2 8 38 126 AND $T=22280 21740 0 0 $X=22290 $Y=21740
X287 3 6 2 11 14 127 AND $T=26680 21740 0 0 $X=26690 $Y=21740
X288 9 6 2 11 33 131 AND $T=31080 21740 0 0 $X=31090 $Y=21740
X289 46 2 6 35 30 31 73 74 225 half_adder $T=50 21780 1 0 $X=50 $Y=17980
X290 50 2 6 26 13 24 102 103 228 half_adder $T=17640 14460 1 0 $X=17640 $Y=10660
X291 22 2 6 25 17 27 129 130 237 half_adder $T=29830 14460 1 0 $X=29830 $Y=10660
X292 43 2 6 33 18 40 133 134 238 half_adder $T=34210 21780 1 0 $X=34210 $Y=17980
X293 30 6 47 2 41 34 44 67 70 71
+ 65 66 68 69 223 224 full_adder1_small $T=22270 7090 1 180 $X=20 $Y=7100
X294 19 6 23 2 42 10 12 60 63 64
+ 58 59 61 62 221 222 full_adder1_small $T=30 -230 0 0 $X=50 $Y=-220
X295 29 6 31 2 44 21 23 53 56 57
+ 51 52 54 55 219 220 full_adder1_small $T=30 7150 1 0 $X=50 $Y=3340
X296 45 6 49 2 39 37 35 86 89 90
+ 84 85 87 88 226 227 full_adder1_small $T=12230 21790 1 0 $X=12250 $Y=17980
X297 38 6 32 2 40 25 39 96 99 100
+ 94 95 97 98 229 230 full_adder1_small $T=17850 14410 0 0 $X=17870 $Y=14420
X298 20 6 21 2 28 15 42 121 124 125
+ 119 120 122 123 235 236 full_adder1_small $T=21990 -230 0 0 $X=22010 $Y=-220
X299 36 6 34 2 24 16 28 114 117 118
+ 112 113 115 116 233 234 full_adder1_small $T=21990 7150 1 0 $X=22010 $Y=3340
X300 48 6 37 2 27 26 41 107 110 111
+ 105 106 108 109 231 232 full_adder1_small $T=21990 7090 0 0 $X=22010 $Y=7100
M0 77 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=11610 $dt=1
M1 76 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=16790 $dt=1
M2 75 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=17.6697 scb=0.0185533 scc=0.000444231 $X=740 $Y=24110 $dt=1
M3 73 46 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=16.2188 scb=0.0173423 scc=0.000698846 $X=750 $Y=18640 $dt=1
M4 58 19 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=2120 $dt=1
M5 51 29 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=4320 $dt=1
M6 44 71 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=1070 $Y=9450 $dt=1
M7 6 70 44 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=1480 $Y=9450 $dt=1
M8 59 23 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=2120 $dt=1
M9 52 31 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=4320 $dt=1
M10 77 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=11600 $dt=1
M11 76 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=16800 $dt=1
M12 75 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1525 scb=0.00906354 scc=0.000187093 $X=1980 $Y=24120 $dt=1
M13 221 23 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=1880 $dt=1
M14 219 31 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=4080 $dt=1
M15 19 77 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=11580 $dt=1
M16 29 76 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=16820 $dt=1
M17 45 75 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=3660 $Y=24140 $dt=1
M18 71 47 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=3910 $Y=9450 $dt=1
M19 60 58 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=1940 $dt=1
M20 53 51 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=4020 $dt=1
M21 6 30 71 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=4320 $Y=9450 $dt=1
M22 60 59 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=1940 $dt=1
M23 53 52 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=4020 $dt=1
M24 80 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=11610 $dt=1
M25 79 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=16790 $dt=1
M26 78 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=5140 $Y=24110 $dt=1
M27 221 19 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=1940 $dt=1
M28 219 29 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=4020 $dt=1
M29 30 35 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=6190 $Y=18700 $dt=1
M30 80 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=11600 $dt=1
M31 79 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=16800 $dt=1
M32 78 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=6380 $Y=24120 $dt=1
M33 70 67 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=6890 $Y=9230 $dt=1
M34 6 41 70 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=7300 $Y=9230 $dt=1
M35 30 46 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=7300 $Y=18660 $dt=1
M36 61 42 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=2120 $dt=1
M37 54 44 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=4320 $dt=1
M38 20 80 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=11580 $dt=1
M39 47 79 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=16820 $dt=1
M40 46 78 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=8060 $Y=24140 $dt=1
M41 74 46 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=8540 $Y=18930 $dt=1
M42 62 60 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=2120 $dt=1
M43 55 53 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=4320 $dt=1
M44 6 41 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=9370 $Y=9260 $dt=1
M45 83 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=11610 $dt=1
M46 82 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=16790 $dt=1
M47 81 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=9540 $Y=24110 $dt=1
M48 74 35 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=9780 $Y=18920 $dt=1
M49 222 60 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=1880 $dt=1
M50 220 53 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=4080 $dt=1
M51 224 69 34 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10330 $Y=9260 $dt=1
M52 83 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=11600 $dt=1
M53 82 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=16800 $dt=1
M54 81 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=10780 $Y=24120 $dt=1
M55 10 61 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=1940 $dt=1
M56 21 54 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=4020 $dt=1
M57 224 68 34 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11290 $Y=9260 $dt=1
M58 31 74 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=11460 $Y=18900 $dt=1
M59 10 62 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=1940 $dt=1
M60 21 55 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=4020 $dt=1
M61 6 67 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=12260 $Y=9200 $dt=1
M62 36 83 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=11580 $dt=1
M63 48 82 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=16820 $dt=1
M64 32 81 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=12460 $Y=24140 $dt=1
M65 222 42 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=1940 $dt=1
M66 220 44 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=4020 $dt=1
M67 84 45 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13020 $Y=18960 $dt=1
M68 6 67 69 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13590 $Y=9440 $dt=1
M69 93 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=11610 $dt=1
M70 92 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=16790 $dt=1
M71 91 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=13940 $Y=24110 $dt=1
M72 85 49 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13980 $Y=18960 $dt=1
M73 6 41 68 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=14550 $Y=9440 $dt=1
M74 63 42 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=1910 $dt=1
M75 56 44 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=4050 $dt=1
M76 93 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=11600 $dt=1
M77 92 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=16800 $dt=1
M78 91 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=15180 $Y=24120 $dt=1
M79 226 49 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=15310 $Y=18720 $dt=1
M80 6 60 63 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=1910 $dt=1
M81 6 53 56 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=4050 $dt=1
M82 6 30 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16210 $Y=9260 $dt=1
M83 86 84 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16280 $Y=18660 $dt=1
M84 50 93 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=11580 $dt=1
M85 22 92 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=16820 $dt=1
M86 49 91 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=16860 $Y=24140 $dt=1
M87 223 66 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17170 $Y=9260 $dt=1
M88 86 85 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17240 $Y=18660 $dt=1
M89 64 19 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=2130 $dt=1
M90 57 29 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=4310 $dt=1
M91 223 65 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18130 $Y=9260 $dt=1
M92 226 45 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18200 $Y=18660 $dt=1
M93 6 23 64 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=2130 $dt=1
M94 6 31 57 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=4310 $dt=1
M95 102 50 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=18340 $Y=11320 $dt=1
M96 104 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=18580 $Y=24110 $dt=1
M97 94 38 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=18640 $Y=16760 $dt=1
M98 6 47 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=19100 $Y=9200 $dt=1
M99 95 32 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19600 $Y=16760 $dt=1
M100 104 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=19820 $Y=24120 $dt=1
M101 87 39 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19860 $Y=18960 $dt=1
M102 6 47 66 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20430 $Y=9440 $dt=1
M103 12 63 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=2130 $dt=1
M104 23 56 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=4310 $dt=1
M105 88 86 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20820 $Y=18960 $dt=1
M106 229 32 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=20930 $Y=16520 $dt=1
M107 6 64 12 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=2130 $dt=1
M108 6 57 23 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=4310 $dt=1
M109 6 30 65 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=21390 $Y=9440 $dt=1
M110 43 104 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=21500 $Y=24140 $dt=1
M111 96 94 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=21900 $Y=16580 $dt=1
M112 227 86 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=22150 $Y=18720 $dt=1
M113 119 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=2120 $dt=1
M114 112 36 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=4320 $dt=1
M115 105 48 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=9440 $dt=1
M116 96 95 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=22860 $Y=16580 $dt=1
M117 126 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=22980 $Y=24110 $dt=1
M118 37 87 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23120 $Y=18660 $dt=1
M119 120 21 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=2120 $dt=1
M120 113 34 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=4320 $dt=1
M121 106 37 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=9440 $dt=1
M122 13 26 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=23780 $Y=11380 $dt=1
M123 229 38 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23820 $Y=16580 $dt=1
M124 37 88 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24080 $Y=18660 $dt=1
M125 126 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=24220 $Y=24120 $dt=1
M126 13 50 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24890 $Y=11340 $dt=1
M127 227 39 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=25040 $Y=18660 $dt=1
M128 235 21 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=1880 $dt=1
M129 233 34 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=4080 $dt=1
M130 231 37 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=9200 $dt=1
M131 97 40 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=25480 $Y=16760 $dt=1
M132 38 126 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=25900 $Y=24140 $dt=1
M133 121 119 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=1940 $dt=1
M134 114 112 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=4020 $dt=1
M135 107 105 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=9260 $dt=1
M136 103 50 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26130 $Y=11610 $dt=1
M137 98 96 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=26440 $Y=16760 $dt=1
M138 121 120 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=1940 $dt=1
M139 114 113 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=4020 $dt=1
M140 107 106 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=9260 $dt=1
M141 89 39 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27110 $Y=18690 $dt=1
M142 103 26 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27370 $Y=11600 $dt=1
M143 127 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=27380 $Y=24110 $dt=1
M144 6 86 89 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27520 $Y=18690 $dt=1
M145 230 96 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=27770 $Y=16520 $dt=1
M146 235 20 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=1940 $dt=1
M147 233 36 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=4020 $dt=1
M148 231 48 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=9260 $dt=1
M149 127 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=28620 $Y=24120 $dt=1
M150 25 97 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28740 $Y=16580 $dt=1
M151 24 103 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=29050 $Y=11580 $dt=1
M152 122 28 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=2120 $dt=1
M153 115 24 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=4320 $dt=1
M154 108 27 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=9440 $dt=1
M155 25 98 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=29700 $Y=16580 $dt=1
M156 90 45 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30090 $Y=18950 $dt=1
M157 14 127 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=30300 $Y=24140 $dt=1
M158 6 49 90 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30500 $Y=18950 $dt=1
M159 129 22 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=30530 $Y=11320 $dt=1
M160 123 121 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=2120 $dt=1
M161 116 114 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=4320 $dt=1
M162 109 107 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=9440 $dt=1
M163 230 40 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=30660 $Y=16580 $dt=1
M164 131 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=31780 $Y=24110 $dt=1
M165 236 121 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=1880 $dt=1
M166 234 114 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=4080 $dt=1
M167 232 107 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=9200 $dt=1
M168 99 40 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=32730 $Y=16550 $dt=1
M169 15 122 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=1940 $dt=1
M170 16 115 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=4020 $dt=1
M171 26 108 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=9260 $dt=1
M172 35 89 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=32930 $Y=18950 $dt=1
M173 131 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=33020 $Y=24120 $dt=1
M174 6 96 99 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=33140 $Y=16550 $dt=1
M175 6 90 35 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=33340 $Y=18950 $dt=1
M176 15 123 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=1940 $dt=1
M177 16 116 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=4020 $dt=1
M178 26 109 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=9260 $dt=1
M179 33 131 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.059 scb=0.0122627 scc=0.000187408 $X=34700 $Y=24140 $dt=1
M180 236 28 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=1940 $dt=1
M181 234 24 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=4020 $dt=1
M182 232 27 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=9260 $dt=1
M183 133 43 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=34910 $Y=18640 $dt=1
M184 100 38 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=35710 $Y=16770 $dt=1
M185 17 25 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=35970 $Y=11380 $dt=1
M186 6 32 100 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=36120 $Y=16770 $dt=1
M187 124 28 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=1910 $dt=1
M188 117 24 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=4050 $dt=1
M189 110 27 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=9230 $dt=1
M190 17 22 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=37080 $Y=11340 $dt=1
M191 6 121 124 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=1910 $dt=1
M192 6 114 117 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=4050 $dt=1
M193 6 107 110 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=9230 $dt=1
M194 130 22 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=38320 $Y=11610 $dt=1
M195 39 99 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=38550 $Y=16770 $dt=1
M196 6 100 39 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=38960 $Y=16770 $dt=1
M197 130 25 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=39560 $Y=11600 $dt=1
M198 125 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=2130 $dt=1
M199 118 36 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=4310 $dt=1
M200 111 48 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=9450 $dt=1
M201 6 21 125 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=2130 $dt=1
M202 6 34 118 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=4310 $dt=1
M203 6 37 111 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=9450 $dt=1
M204 18 33 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.2705 scb=0.0126902 scc=0.000796523 $X=40350 $Y=18700 $dt=1
M205 27 130 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=41240 $Y=11580 $dt=1
M206 18 43 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=41460 $Y=18660 $dt=1
M207 42 124 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=2130 $dt=1
M208 28 117 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=4310 $dt=1
M209 41 110 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=42690 $Y=9450 $dt=1
M210 134 43 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42700 $Y=18930 $dt=1
M211 6 125 42 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=2130 $dt=1
M212 6 118 28 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=4310 $dt=1
M213 6 111 41 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=43100 $Y=9450 $dt=1
M214 134 33 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43940 $Y=18920 $dt=1
M215 40 134 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=45620 $Y=18900 $dt=1
.ends multiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_31                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_31 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_31

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_32                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_32 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_32

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_43                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_43 1 2 3 5 6 8
** N=14 EP=6 FDC=4
M0 8 6 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=810 $Y=710 $dt=0
M1 5 3 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=4640 $Y=580 $dt=0
M2 8 6 1 1 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=810 $Y=2230 $dt=1
M3 5 3 1 1 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.2373 scb=0.0194294 scc=0.00149528 $X=4640 $Y=1900 $dt=1
.ends cellTmpl_CDNS_43

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_44                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_44 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_44

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_45                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_45 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_45

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=12
X0 7 M3_M2_CDNS_8 $T=250 -3000 0 0 $X=170 $Y=-3250
X1 7 M3_M2_CDNS_8 $T=960 -2040 0 0 $X=880 $Y=-2290
X2 7 M3_M2_CDNS_8 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X3 7 M2_M1_CDNS_9 $T=960 -2040 0 0 $X=880 $Y=-2290
X4 1 M1_PO_CDNS_13 $T=1300 -3500 0 0 $X=1200 $Y=-3750
X5 1 M1_PO_CDNS_13 $T=2660 -4240 0 0 $X=2560 $Y=-4490
X6 1 M1_PO_CDNS_14 $T=680 -3550 0 0 $X=580 $Y=-3670
X7 2 M1_PO_CDNS_14 $T=1300 -2090 0 0 $X=1200 $Y=-2210
X8 5 M1_PO_CDNS_14 $T=4040 -3180 0 0 $X=3940 $Y=-3300
X9 8 M1_PO_CDNS_14 $T=4300 -3670 0 90 $X=4180 $Y=-3770
X10 1 M2_M1_CDNS_15 $T=1300 -3500 0 0 $X=1220 $Y=-3750
X11 1 M2_M1_CDNS_15 $T=2660 -4240 0 0 $X=2580 $Y=-4490
X12 7 M2_M1_CDNS_16 $T=250 -3000 0 0 $X=170 $Y=-3250
X13 7 M2_M1_CDNS_16 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X14 7 M1_PO_CDNS_17 $T=250 -3000 0 0 $X=150 $Y=-3250
X15 7 M1_PO_CDNS_17 $T=2620 -2730 0 0 $X=2520 $Y=-2980
X16 4 7 9 4 nmos1v_CDNS_31 $T=1990 -4420 0 0 $X=1790 $Y=-4620
X17 8 5 10 4 nmos1v_CDNS_31 $T=3370 -4430 0 0 $X=3170 $Y=-4630
X18 8 2 9 4 nmos1v_CDNS_32 $T=1780 -4420 0 0 $X=1360 $Y=-4620
X19 4 1 10 4 nmos1v_CDNS_32 $T=3160 -4430 0 0 $X=2740 $Y=-4630
X20 3 4 8 6 1 7 cellTmpl_CDNS_43 $T=-60 -5080 0 0 $X=-180 $Y=-5220
X21 3 1 11 4 3 pmos1v_CDNS_44 $T=1990 -3120 0 0 $X=1790 $Y=-3320
X22 8 5 12 4 3 pmos1v_CDNS_44 $T=3370 -3190 0 0 $X=3170 $Y=-3390
X23 8 2 11 4 3 pmos1v_CDNS_45 $T=1780 -3120 0 0 $X=1360 $Y=-3320
X24 3 7 12 4 3 pmos1v_CDNS_45 $T=3160 -3190 0 0 $X=2740 $Y=-3390
M0 9 2 8 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1780 $Y=-4420 $dt=0
M1 4 7 9 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1990 $Y=-4420 $dt=0
M2 10 1 4 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3160 $Y=-4430 $dt=0
M3 8 5 10 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3370 $Y=-4430 $dt=0
M4 11 2 8 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1780 $Y=-3120 $dt=1
M5 3 1 11 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1990 $Y=-3120 $dt=1
M6 12 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3160 $Y=-3190 $dt=1
M7 8 5 12 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3370 $Y=-3190 $dt=1
.ends MUX_2to1___2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FA_4bit                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FA_4bit 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19
** N=83 EP=19 FDC=144
X0 5 M2_M1_CDNS_1 $T=-80 3540 0 0 $X=-160 $Y=3410
X1 5 M2_M1_CDNS_1 $T=-80 10890 0 0 $X=-160 $Y=10760
X2 17 M2_M1_CDNS_1 $T=21770 2020 0 0 $X=21690 $Y=1890
X3 18 M2_M1_CDNS_1 $T=21770 5100 0 0 $X=21690 $Y=4970
X4 18 M3_M2_CDNS_2 $T=21980 9220 0 0 $X=21900 $Y=9090
X5 17 M4_M3_CDNS_3 $T=14030 6120 0 0 $X=13950 $Y=5870
X6 19 M4_M3_CDNS_3 $T=16960 11880 0 0 $X=16880 $Y=11630
X7 17 M4_M3_CDNS_3 $T=19730 4760 0 0 $X=19650 $Y=4510
X8 19 M4_M3_CDNS_3 $T=22610 11350 0 0 $X=22530 $Y=11100
X9 17 M3_M2_CDNS_6 $T=14030 6120 0 0 $X=13950 $Y=5870
X10 19 M3_M2_CDNS_6 $T=16960 11880 0 0 $X=16880 $Y=11630
X11 19 M3_M2_CDNS_6 $T=22610 11350 0 0 $X=22530 $Y=11100
X12 17 M3_M2_CDNS_7 $T=19730 4760 0 0 $X=19650 $Y=4510
X13 18 M3_M2_CDNS_8 $T=18840 8310 0 0 $X=18760 $Y=8060
X14 17 M2_M1_CDNS_16 $T=14030 6120 0 0 $X=13950 $Y=5870
X15 19 M2_M1_CDNS_16 $T=16960 11880 0 0 $X=16880 $Y=11630
X16 18 M2_M1_CDNS_16 $T=18840 8310 0 0 $X=18760 $Y=8060
X17 19 M2_M1_CDNS_16 $T=22610 11350 0 0 $X=22530 $Y=11100
X18 17 M1_PO_CDNS_17 $T=14030 6120 0 0 $X=13930 $Y=5870
X19 19 M1_PO_CDNS_17 $T=16960 11880 0 0 $X=16860 $Y=11630
X20 18 M1_PO_CDNS_17 $T=18840 8310 0 0 $X=18740 $Y=8060
X21 6 5 1 7 11 12 17 43 46 47
+ 41 42 44 45 82 83 full_adder1_small $T=-90 -130 0 0 $X=-70 $Y=-120
X22 8 5 2 7 17 13 18 36 39 40
+ 34 35 37 38 80 81 full_adder1_small $T=-90 7250 1 0 $X=-70 $Y=3440
X23 9 5 3 7 18 14 19 29 32 33
+ 27 28 30 31 78 79 full_adder1_small $T=-90 7190 0 0 $X=-70 $Y=7200
X24 10 5 4 7 19 15 16 22 25 26
+ 20 21 23 24 76 77 full_adder1_small $T=-90 14570 1 0 $X=-70 $Y=10760
M0 41 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=2220 $dt=1
M1 34 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=4420 $dt=1
M2 27 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=9540 $dt=1
M3 20 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=11740 $dt=1
M4 42 1 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=2220 $dt=1
M5 35 2 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=4420 $dt=1
M6 28 3 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=9540 $dt=1
M7 21 4 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=11740 $dt=1
M8 82 1 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=1980 $dt=1
M9 80 2 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=4180 $dt=1
M10 78 3 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=9300 $dt=1
M11 76 4 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=11500 $dt=1
M12 43 41 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=2040 $dt=1
M13 36 34 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=4120 $dt=1
M14 29 27 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=9360 $dt=1
M15 22 20 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=11440 $dt=1
M16 43 42 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=2040 $dt=1
M17 36 35 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=4120 $dt=1
M18 29 28 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=9360 $dt=1
M19 22 21 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=11440 $dt=1
M20 82 6 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=2040 $dt=1
M21 80 8 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=4120 $dt=1
M22 78 9 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=9360 $dt=1
M23 76 10 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=11440 $dt=1
M24 44 11 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=2220 $dt=1
M25 37 17 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=4420 $dt=1
M26 30 18 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=9540 $dt=1
M27 23 19 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=11740 $dt=1
M28 45 43 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=2220 $dt=1
M29 38 36 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=4420 $dt=1
M30 31 29 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=9540 $dt=1
M31 24 22 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=11740 $dt=1
M32 83 43 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=1980 $dt=1
M33 81 36 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=4180 $dt=1
M34 79 29 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=9300 $dt=1
M35 77 22 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=11500 $dt=1
M36 12 44 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=2040 $dt=1
M37 13 37 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=4120 $dt=1
M38 14 30 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=9360 $dt=1
M39 15 23 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=11440 $dt=1
M40 12 45 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=2040 $dt=1
M41 13 38 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=4120 $dt=1
M42 14 31 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=9360 $dt=1
M43 15 24 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=11440 $dt=1
M44 83 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=2040 $dt=1
M45 81 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=4120 $dt=1
M46 79 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=9360 $dt=1
M47 77 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=11440 $dt=1
M48 46 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=2010 $dt=1
M49 39 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=4150 $dt=1
M50 32 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=9330 $dt=1
M51 25 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=11470 $dt=1
M52 5 43 46 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=2010 $dt=1
M53 5 36 39 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=4150 $dt=1
M54 5 29 32 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=9330 $dt=1
M55 5 22 25 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=11470 $dt=1
M56 47 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=2230 $dt=1
M57 40 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=4410 $dt=1
M58 33 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=9550 $dt=1
M59 26 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=11730 $dt=1
M60 5 1 47 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=2230 $dt=1
M61 5 2 40 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=4410 $dt=1
M62 5 3 33 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=9550 $dt=1
M63 5 4 26 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=11730 $dt=1
M64 17 46 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=2230 $dt=1
M65 18 39 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=4410 $dt=1
M66 19 32 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=9550 $dt=1
M67 16 25 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=11730 $dt=1
M68 5 47 17 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=2230 $dt=1
M69 5 40 18 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=4410 $dt=1
M70 5 33 19 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=9550 $dt=1
M71 5 26 16 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=11730 $dt=1
.ends FA_4bit

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small 1 2 3 4
** N=4 EP=4 FDC=2
X0 1 M1_PO_CDNS_14 $T=950 1780 0 90 $X=830 $Y=1680
X1 2 3 cellTmpl_CDNS_18 $T=120 140 0 0 $X=0 $Y=0
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7353 scb=0.0117274 scc=0.000445561 $X=1070 $Y=980 $dt=0
M1 4 1 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8675 scb=0.0146094 scc=0.000688105 $X=1070 $Y=2220 $dt=1
.ends INV_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 10badder                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 10badder 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59
** N=267 EP=59 FDC=516
X0 3 M2_M1_CDNS_1 $T=50480 50560 0 0 $X=50400 $Y=50430
X1 3 M2_M1_CDNS_1 $T=51590 45750 0 90 $X=51460 $Y=45670
X2 35 M2_M1_CDNS_1 $T=53210 27000 0 0 $X=53130 $Y=26870
X3 36 M2_M1_CDNS_1 $T=53210 41640 0 0 $X=53130 $Y=41510
X4 37 M2_M1_CDNS_1 $T=53230 23140 0 0 $X=53150 $Y=23010
X5 38 M2_M1_CDNS_1 $T=53230 37780 0 0 $X=53150 $Y=37650
X6 3 M2_M1_CDNS_1 $T=62920 24380 0 0 $X=62840 $Y=24250
X7 3 M2_M1_CDNS_1 $T=62920 39020 0 0 $X=62840 $Y=38890
X8 3 M2_M1_CDNS_1 $T=62930 31710 0 0 $X=62850 $Y=31580
X9 3 M2_M1_CDNS_1 $T=62930 46350 0 0 $X=62850 $Y=46220
X10 35 M3_M2_CDNS_2 $T=50730 34460 0 0 $X=50650 $Y=34330
X11 36 M3_M2_CDNS_2 $T=50800 49100 0 0 $X=50720 $Y=48970
X12 2 M3_M2_CDNS_2 $T=51610 22610 0 0 $X=51530 $Y=22480
X13 39 M4_M3_CDNS_3 $T=51080 34160 0 0 $X=51000 $Y=33910
X14 40 M4_M3_CDNS_3 $T=56340 32800 0 0 $X=56260 $Y=32550
X15 41 M4_M3_CDNS_3 $T=56340 47440 0 0 $X=56260 $Y=47190
X16 42 M4_M3_CDNS_3 $T=57240 50840 0 0 $X=57160 $Y=50590
X17 43 M4_M3_CDNS_3 $T=72650 52420 0 90 $X=72400 $Y=52340
X18 39 M4_M3_CDNS_3 $T=78550 36430 0 0 $X=78470 $Y=36180
X19 43 M4_M3_CDNS_3 $T=79400 52420 0 90 $X=79150 $Y=52340
X20 40 M4_M3_CDNS_3 $T=86760 34460 0 0 $X=86680 $Y=34210
X21 41 M4_M3_CDNS_3 $T=86760 49100 0 0 $X=86680 $Y=48850
X22 39 M4_M3_CDNS_5 $T=51140 36930 0 0 $X=51060 $Y=36800
X23 39 M3_M2_CDNS_6 $T=51080 34160 0 0 $X=51000 $Y=33910
X24 40 M3_M2_CDNS_6 $T=56340 32800 0 0 $X=56260 $Y=32550
X25 41 M3_M2_CDNS_6 $T=56340 47440 0 0 $X=56260 $Y=47190
X26 42 M3_M2_CDNS_6 $T=57240 50840 0 0 $X=57160 $Y=50590
X27 43 M3_M2_CDNS_6 $T=72650 52420 0 90 $X=72400 $Y=52340
X28 39 M3_M2_CDNS_6 $T=78550 36430 0 0 $X=78470 $Y=36180
X29 43 M3_M2_CDNS_6 $T=79400 52420 0 90 $X=79150 $Y=52340
X30 40 M3_M2_CDNS_6 $T=86760 34460 0 0 $X=86680 $Y=34210
X31 41 M3_M2_CDNS_6 $T=86760 49100 0 0 $X=86680 $Y=48850
X32 2 M3_M2_CDNS_8 $T=52330 32180 0 90 $X=52080 $Y=32100
X33 39 M3_M2_CDNS_8 $T=52330 46820 0 90 $X=52080 $Y=46740
X34 44 M3_M2_CDNS_8 $T=53480 29020 0 0 $X=53400 $Y=28770
X35 45 M3_M2_CDNS_8 $T=53480 43660 0 0 $X=53400 $Y=43410
X36 46 M3_M2_CDNS_8 $T=54270 29810 0 90 $X=54020 $Y=29730
X37 47 M3_M2_CDNS_8 $T=54270 44450 0 90 $X=54020 $Y=44370
X38 44 M3_M2_CDNS_8 $T=55540 26280 0 0 $X=55460 $Y=26030
X39 45 M3_M2_CDNS_8 $T=55540 40920 0 0 $X=55460 $Y=40670
X40 48 M3_M2_CDNS_8 $T=55730 21200 0 90 $X=55480 $Y=21120
X41 49 M3_M2_CDNS_8 $T=55730 35840 0 90 $X=55480 $Y=35760
X42 50 M3_M2_CDNS_8 $T=56210 23810 0 90 $X=55960 $Y=23730
X43 51 M3_M2_CDNS_8 $T=56210 38450 0 90 $X=55960 $Y=38370
X44 52 M3_M2_CDNS_8 $T=56050 31070 0 0 $X=55970 $Y=30820
X45 53 M3_M2_CDNS_8 $T=56050 45710 0 0 $X=55970 $Y=45460
X46 35 M3_M2_CDNS_8 $T=56240 34220 0 0 $X=56160 $Y=33970
X47 36 M3_M2_CDNS_8 $T=56240 48860 0 0 $X=56160 $Y=48610
X48 13 M3_M2_CDNS_8 $T=57660 26200 0 90 $X=57410 $Y=26120
X49 11 M3_M2_CDNS_8 $T=57660 33520 0 90 $X=57410 $Y=33440
X50 10 M3_M2_CDNS_8 $T=57660 40840 0 90 $X=57410 $Y=40760
X51 8 M3_M2_CDNS_8 $T=57660 48160 0 90 $X=57410 $Y=48080
X52 7 M3_M2_CDNS_8 $T=57670 22770 0 90 $X=57420 $Y=22690
X53 12 M3_M2_CDNS_8 $T=57670 30070 0 90 $X=57420 $Y=29990
X54 6 M3_M2_CDNS_8 $T=57670 37410 0 90 $X=57420 $Y=37330
X55 9 M3_M2_CDNS_8 $T=57670 44710 0 90 $X=57420 $Y=44630
X56 52 M3_M2_CDNS_8 $T=62950 31240 0 90 $X=62700 $Y=31160
X57 53 M3_M2_CDNS_8 $T=62950 45880 0 90 $X=62700 $Y=45800
X58 50 M3_M2_CDNS_8 $T=63400 23460 0 0 $X=63320 $Y=23210
X59 51 M3_M2_CDNS_8 $T=63400 38100 0 0 $X=63320 $Y=37850
X60 48 M3_M2_CDNS_8 $T=63720 21760 0 0 $X=63640 $Y=21510
X61 49 M3_M2_CDNS_8 $T=63720 36400 0 0 $X=63640 $Y=36150
X62 46 M3_M2_CDNS_8 $T=63820 29420 0 0 $X=63740 $Y=29170
X63 47 M3_M2_CDNS_8 $T=63820 44060 0 0 $X=63740 $Y=43810
X64 44 M2_M1_CDNS_9 $T=53480 29020 0 0 $X=53400 $Y=28770
X65 45 M2_M1_CDNS_9 $T=53480 43660 0 0 $X=53400 $Y=43410
X66 35 M2_M1_CDNS_9 $T=56240 34220 0 0 $X=56160 $Y=33970
X67 36 M2_M1_CDNS_9 $T=56240 48860 0 0 $X=56160 $Y=48610
X68 52 M2_M1_CDNS_9 $T=62950 31240 0 90 $X=62700 $Y=31160
X69 53 M2_M1_CDNS_9 $T=62950 45880 0 90 $X=62700 $Y=45800
X70 50 M2_M1_CDNS_9 $T=63400 23460 0 0 $X=63320 $Y=23210
X71 51 M2_M1_CDNS_9 $T=63400 38100 0 0 $X=63320 $Y=37850
X72 48 M2_M1_CDNS_9 $T=63720 21760 0 0 $X=63640 $Y=21510
X73 49 M2_M1_CDNS_9 $T=63720 36400 0 0 $X=63640 $Y=36150
X74 46 M2_M1_CDNS_9 $T=63820 29420 0 0 $X=63740 $Y=29170
X75 47 M2_M1_CDNS_9 $T=63820 44060 0 0 $X=63740 $Y=43810
X76 37 M1_PO_CDNS_13 $T=53520 24980 0 90 $X=53270 $Y=24880
X77 38 M1_PO_CDNS_13 $T=53520 39620 0 90 $X=53270 $Y=39520
X78 14 M1_PO_CDNS_13 $T=64110 23330 0 0 $X=64010 $Y=23080
X79 18 M1_PO_CDNS_13 $T=64110 37970 0 0 $X=64010 $Y=37720
X80 14 M1_PO_CDNS_13 $T=65950 23850 0 90 $X=65700 $Y=23750
X81 18 M1_PO_CDNS_13 $T=65950 38490 0 90 $X=65700 $Y=38390
X82 2 M1_PO_CDNS_13 $T=78510 22370 0 0 $X=78410 $Y=22120
X83 54 M1_PO_CDNS_14 $T=53270 31100 0 0 $X=53170 $Y=30980
X84 55 M1_PO_CDNS_14 $T=53270 45740 0 0 $X=53170 $Y=45620
X85 56 M1_PO_CDNS_14 $T=53550 23450 0 0 $X=53450 $Y=23330
X86 57 M1_PO_CDNS_14 $T=53550 38090 0 0 $X=53450 $Y=37970
X87 58 M1_PO_CDNS_14 $T=53840 25910 0 0 $X=53740 $Y=25790
X88 59 M1_PO_CDNS_14 $T=53840 40550 0 0 $X=53740 $Y=40430
X89 37 M2_M1_CDNS_15 $T=53520 24980 0 90 $X=53270 $Y=24900
X90 38 M2_M1_CDNS_15 $T=53520 39620 0 90 $X=53270 $Y=39540
X91 14 M2_M1_CDNS_15 $T=64110 23330 0 0 $X=64030 $Y=23080
X92 18 M2_M1_CDNS_15 $T=64110 37970 0 0 $X=64030 $Y=37720
X93 14 M2_M1_CDNS_15 $T=65950 23850 0 90 $X=65700 $Y=23770
X94 18 M2_M1_CDNS_15 $T=65950 38490 0 90 $X=65700 $Y=38410
X95 2 M2_M1_CDNS_15 $T=78510 22370 0 0 $X=78430 $Y=22120
X96 39 M2_M1_CDNS_16 $T=51080 34160 0 0 $X=51000 $Y=33910
X97 2 M2_M1_CDNS_16 $T=52330 32180 0 90 $X=52080 $Y=32100
X98 39 M2_M1_CDNS_16 $T=52330 46820 0 90 $X=52080 $Y=46740
X99 46 M2_M1_CDNS_16 $T=54270 29810 0 90 $X=54020 $Y=29730
X100 47 M2_M1_CDNS_16 $T=54270 44450 0 90 $X=54020 $Y=44370
X101 44 M2_M1_CDNS_16 $T=55540 26280 0 0 $X=55460 $Y=26030
X102 45 M2_M1_CDNS_16 $T=55540 40920 0 0 $X=55460 $Y=40670
X103 48 M2_M1_CDNS_16 $T=55730 21200 0 90 $X=55480 $Y=21120
X104 49 M2_M1_CDNS_16 $T=55730 35840 0 90 $X=55480 $Y=35760
X105 50 M2_M1_CDNS_16 $T=56210 23810 0 90 $X=55960 $Y=23730
X106 51 M2_M1_CDNS_16 $T=56210 38450 0 90 $X=55960 $Y=38370
X107 52 M2_M1_CDNS_16 $T=56050 31070 0 0 $X=55970 $Y=30820
X108 53 M2_M1_CDNS_16 $T=56050 45710 0 0 $X=55970 $Y=45460
X109 40 M2_M1_CDNS_16 $T=56340 32800 0 0 $X=56260 $Y=32550
X110 41 M2_M1_CDNS_16 $T=56340 47440 0 0 $X=56260 $Y=47190
X111 42 M2_M1_CDNS_16 $T=57240 50840 0 0 $X=57160 $Y=50590
X112 13 M2_M1_CDNS_16 $T=57660 26200 0 90 $X=57410 $Y=26120
X113 11 M2_M1_CDNS_16 $T=57660 33520 0 90 $X=57410 $Y=33440
X114 10 M2_M1_CDNS_16 $T=57660 40840 0 90 $X=57410 $Y=40760
X115 8 M2_M1_CDNS_16 $T=57660 48160 0 90 $X=57410 $Y=48080
X116 7 M2_M1_CDNS_16 $T=57670 22770 0 90 $X=57420 $Y=22690
X117 12 M2_M1_CDNS_16 $T=57670 30070 0 90 $X=57420 $Y=29990
X118 6 M2_M1_CDNS_16 $T=57670 37410 0 90 $X=57420 $Y=37330
X119 9 M2_M1_CDNS_16 $T=57670 44710 0 90 $X=57420 $Y=44630
X120 43 M2_M1_CDNS_16 $T=72650 52420 0 90 $X=72400 $Y=52340
X121 39 M2_M1_CDNS_16 $T=78550 36430 0 0 $X=78470 $Y=36180
X122 43 M2_M1_CDNS_16 $T=79400 52420 0 90 $X=79150 $Y=52340
X123 40 M2_M1_CDNS_16 $T=86760 34460 0 0 $X=86680 $Y=34210
X124 41 M2_M1_CDNS_16 $T=86760 49100 0 0 $X=86680 $Y=48850
X125 2 M1_PO_CDNS_17 $T=52330 32180 0 90 $X=52080 $Y=32080
X126 39 M1_PO_CDNS_17 $T=52330 46820 0 90 $X=52080 $Y=46720
X127 46 M1_PO_CDNS_17 $T=54270 29810 0 90 $X=54020 $Y=29710
X128 47 M1_PO_CDNS_17 $T=54270 44450 0 90 $X=54020 $Y=44350
X129 44 M1_PO_CDNS_17 $T=55540 26280 0 0 $X=55440 $Y=26030
X130 45 M1_PO_CDNS_17 $T=55540 40920 0 0 $X=55440 $Y=40670
X131 48 M1_PO_CDNS_17 $T=55730 21200 0 90 $X=55480 $Y=21100
X132 49 M1_PO_CDNS_17 $T=55730 35840 0 90 $X=55480 $Y=35740
X133 52 M1_PO_CDNS_17 $T=56050 31070 0 0 $X=55950 $Y=30820
X134 53 M1_PO_CDNS_17 $T=56050 45710 0 0 $X=55950 $Y=45460
X135 50 M1_PO_CDNS_17 $T=56210 23810 0 90 $X=55960 $Y=23710
X136 51 M1_PO_CDNS_17 $T=56210 38450 0 90 $X=55960 $Y=38350
X137 40 M1_PO_CDNS_17 $T=56340 32800 0 0 $X=56240 $Y=32550
X138 41 M1_PO_CDNS_17 $T=56340 47440 0 0 $X=56240 $Y=47190
X139 13 M1_PO_CDNS_17 $T=57660 26200 0 90 $X=57410 $Y=26100
X140 11 M1_PO_CDNS_17 $T=57660 33520 0 90 $X=57410 $Y=33420
X141 10 M1_PO_CDNS_17 $T=57660 40840 0 90 $X=57410 $Y=40740
X142 8 M1_PO_CDNS_17 $T=57660 48160 0 90 $X=57410 $Y=48060
X143 7 M1_PO_CDNS_17 $T=57670 22770 0 90 $X=57420 $Y=22670
X144 12 M1_PO_CDNS_17 $T=57670 30070 0 90 $X=57420 $Y=29970
X145 6 M1_PO_CDNS_17 $T=57670 37410 0 90 $X=57420 $Y=37310
X146 9 M1_PO_CDNS_17 $T=57670 44710 0 90 $X=57420 $Y=44610
X147 39 M1_PO_CDNS_17 $T=78550 36430 0 0 $X=78450 $Y=36180
X148 3 4 48 56 50 172 NAND_1X_small $T=53960 20720 0 0 $X=53530 $Y=20700
X149 3 4 44 58 37 171 NAND_1X_small $T=55940 28040 0 180 $X=53530 $Y=24260
X150 3 4 46 54 52 170 NAND_1X_small $T=53960 28040 0 0 $X=53530 $Y=28020
X151 3 4 49 57 51 169 NAND_1X_small $T=53960 35360 0 0 $X=53530 $Y=35340
X152 3 4 45 59 38 168 NAND_1X_small $T=55940 42680 0 180 $X=53530 $Y=38900
X153 3 4 47 55 53 167 NAND_1X_small $T=53960 42680 0 0 $X=53530 $Y=42660
X154 3 4 14 7 50 85 86 187 265 188 XOR1 $T=56070 20720 0 0 $X=56130 $Y=20700
X155 3 4 15 13 48 83 84 185 264 186 XOR1 $T=56070 28040 1 0 $X=56130 $Y=24260
X156 3 4 16 12 52 81 82 183 263 184 XOR1 $T=56070 28040 0 0 $X=56130 $Y=28020
X157 3 4 17 11 46 79 80 181 262 182 XOR1 $T=56070 35360 1 0 $X=56130 $Y=31580
X158 3 4 18 6 51 77 78 179 261 180 XOR1 $T=56070 35360 0 0 $X=56130 $Y=35340
X159 3 4 19 10 49 75 76 177 260 178 XOR1 $T=56070 42680 1 0 $X=56130 $Y=38900
X160 3 4 20 9 53 73 74 175 259 176 XOR1 $T=56070 42680 0 0 $X=56130 $Y=42660
X161 3 4 21 8 47 71 72 173 258 174 XOR1 $T=56070 50000 1 0 $X=56130 $Y=46220
X162 5 3 1 4 42 22 43 66 69 70
+ 64 65 67 68 256 257 full_adder1_small $T=50650 49970 0 0 $X=50670 $Y=49980
X163 24 3 23 4 43 33 34 151 154 155
+ 149 150 152 153 266 267 full_adder1_small $T=72610 49970 0 0 $X=72630 $Y=49980
X164 35 40 3 4 2 39 62 63 158 159
+ 254 255 MUX_2to1___2X $T=56190 30160 0 180 $X=50640 $Y=31580
X165 36 41 3 4 39 42 60 61 156 157
+ 252 253 MUX_2to1___2X $T=56190 44800 0 180 $X=50640 $Y=46220
X166 14 13 12 11 3 7 4 15 16 17
+ 2 25 28 27 26 40 138 140 139 FA_4bit $T=64900 20820 0 0 $X=64250 $Y=20700
X167 18 10 9 8 3 6 4 19 20 21
+ 39 32 31 30 29 41 107 109 108 FA_4bit $T=64900 35460 0 0 $X=64250 $Y=35340
X168 56 3 4 37 INV_1X_small $T=51530 20700 0 0 $X=51530 $Y=20700
X169 58 3 4 35 INV_1X_small $T=51530 28060 1 0 $X=51530 $Y=24260
X170 54 3 4 44 INV_1X_small $T=51530 28020 0 0 $X=51530 $Y=28020
X171 57 3 4 38 INV_1X_small $T=51530 35340 0 0 $X=51530 $Y=35340
X172 59 3 4 36 INV_1X_small $T=51530 42700 1 0 $X=51530 $Y=38900
X173 55 3 4 45 INV_1X_small $T=51530 42660 0 0 $X=51530 $Y=42660
M0 64 5 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6612 scb=0.0167915 scc=0.000377457 $X=51440 $Y=52320 $dt=1
M1 65 1 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.8911 scb=0.00996238 scc=0.000256798 $X=52400 $Y=52320 $dt=1
M2 256 1 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=53730 $Y=52080 $dt=1
M3 58 37 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=25230 $dt=1
M4 59 38 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=39870 $dt=1
M5 66 64 256 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=54700 $Y=52140 $dt=1
M6 56 48 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=23050 $dt=1
M7 54 46 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=30370 $dt=1
M8 57 49 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=37690 $dt=1
M9 55 47 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=45010 $dt=1
M10 3 44 58 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=25230 $dt=1
M11 3 45 59 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=39870 $dt=1
M12 3 50 56 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=23050 $dt=1
M13 3 52 54 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=30370 $dt=1
M14 3 51 57 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=37690 $dt=1
M15 3 53 55 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=45010 $dt=1
M16 66 65 256 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=55660 $Y=52140 $dt=1
M17 256 5 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=56620 $Y=52140 $dt=1
M18 85 14 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=23040 $dt=1
M19 83 15 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=25240 $dt=1
M20 81 16 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=30360 $dt=1
M21 79 17 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=32560 $dt=1
M22 77 18 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=37680 $dt=1
M23 75 19 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=39880 $dt=1
M24 73 20 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=45000 $dt=1
M25 71 21 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=47200 $dt=1
M26 86 7 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=23040 $dt=1
M27 84 13 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=25240 $dt=1
M28 82 12 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=30360 $dt=1
M29 80 11 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=32560 $dt=1
M30 78 6 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=37680 $dt=1
M31 76 10 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=39880 $dt=1
M32 74 9 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=45000 $dt=1
M33 72 8 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=47200 $dt=1
M34 67 42 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=58280 $Y=52320 $dt=1
M35 265 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=22800 $dt=1
M36 264 13 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=25000 $dt=1
M37 263 12 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=30120 $dt=1
M38 262 11 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=32320 $dt=1
M39 261 6 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=37440 $dt=1
M40 260 10 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=39640 $dt=1
M41 259 9 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=44760 $dt=1
M42 258 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=46960 $dt=1
M43 68 66 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=59240 $Y=52320 $dt=1
M44 50 85 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=22860 $dt=1
M45 48 83 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=24940 $dt=1
M46 52 81 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=30180 $dt=1
M47 46 79 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=32260 $dt=1
M48 51 77 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=37500 $dt=1
M49 49 75 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=39580 $dt=1
M50 53 73 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=44820 $dt=1
M51 47 71 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=46900 $dt=1
M52 257 66 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60570 $Y=52080 $dt=1
M53 50 86 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=22860 $dt=1
M54 48 84 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=24940 $dt=1
M55 52 82 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=30180 $dt=1
M56 46 80 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=32260 $dt=1
M57 51 78 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=37500 $dt=1
M58 49 76 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=39580 $dt=1
M59 53 74 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=44820 $dt=1
M60 47 72 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=46900 $dt=1
M61 22 67 257 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=61540 $Y=52140 $dt=1
M62 265 14 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=22860 $dt=1
M63 264 15 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=24940 $dt=1
M64 263 16 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=30180 $dt=1
M65 262 17 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=32260 $dt=1
M66 261 18 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=37500 $dt=1
M67 260 19 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=39580 $dt=1
M68 259 20 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=44820 $dt=1
M69 258 21 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=46900 $dt=1
M70 22 68 257 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=62500 $Y=52140 $dt=1
M71 257 42 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=63460 $Y=52140 $dt=1
M72 69 42 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65530 $Y=52110 $dt=1
M73 3 66 69 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=65940 $Y=52110 $dt=1
M74 70 5 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68510 $Y=52330 $dt=1
M75 3 1 70 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=68920 $Y=52330 $dt=1
M76 43 69 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71350 $Y=52330 $dt=1
M77 3 70 43 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=71760 $Y=52330 $dt=1
M78 149 24 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=73400 $Y=52320 $dt=1
M79 150 23 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=74360 $Y=52320 $dt=1
M80 266 23 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=75690 $Y=52080 $dt=1
M81 151 149 266 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=76660 $Y=52140 $dt=1
M82 151 150 266 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=77620 $Y=52140 $dt=1
M83 266 24 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=78580 $Y=52140 $dt=1
M84 152 43 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=80240 $Y=52320 $dt=1
M85 153 151 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=81200 $Y=52320 $dt=1
M86 267 151 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=82530 $Y=52080 $dt=1
M87 33 152 267 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=83500 $Y=52140 $dt=1
M88 33 153 267 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=84460 $Y=52140 $dt=1
M89 267 43 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=85420 $Y=52140 $dt=1
M90 154 43 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87490 $Y=52110 $dt=1
M91 3 151 154 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=87900 $Y=52110 $dt=1
M92 155 24 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90470 $Y=52330 $dt=1
M93 3 23 155 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=90880 $Y=52330 $dt=1
M94 34 154 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=93310 $Y=52330 $dt=1
M95 3 155 34 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=93720 $Y=52330 $dt=1
.ends 10badder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_46                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_46 1 2 3 5
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=660 $Y=760 $dt=0
.ends cellTmpl_CDNS_46

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 1 M1_PO_CDNS_14 $T=700 2040 0 90 $X=580 $Y=1940
X1 2 3 1 4 cellTmpl_CDNS_46 $T=120 140 0 0 $X=0 $Y=0
.ends INV_1X_small_layout

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_14 $T=640 1830 0 90 $X=520 $Y=1730
X1 6 M1_PO_CDNS_14 $T=1940 640 0 0 $X=1840 $Y=520
X2 3 1 6 3 nmos1v_CDNS_19 $T=710 860 0 0 $X=290 $Y=660
X3 4 6 5 3 nmos1v_CDNS_19 $T=1890 860 0 0 $X=1470 $Y=660
X4 2 3 cellTmpl_CDNS_21 $T=120 140 0 0 $X=0 $Y=0
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=710 $Y=860 $dt=0
M1 5 6 4 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1890 $Y=860 $dt=0
.ends ph1p3_clk_part

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_48                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_48 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_48

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_MSDFF                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_MSDFF 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17
*.DEVICECLIMB
** N=18 EP=17 FDC=15
X0 2 M2_M1_CDNS_1 $T=430 2010 0 0 $X=350 $Y=1880
X1 7 M2_M1_CDNS_1 $T=1110 -1470 0 0 $X=1030 $Y=-1600
X2 2 M2_M1_CDNS_1 $T=2790 -1820 0 0 $X=2710 $Y=-1950
X3 8 M2_M1_CDNS_1 $T=4150 -1460 0 0 $X=4070 $Y=-1590
X4 6 M2_M1_CDNS_1 $T=5200 -2030 0 0 $X=5120 $Y=-2160
X5 7 M2_M1_CDNS_1 $T=5310 1560 0 90 $X=5180 $Y=1480
X6 8 M2_M1_CDNS_1 $T=5670 -1460 0 90 $X=5540 $Y=-1540
X7 9 M2_M1_CDNS_1 $T=6280 1490 0 0 $X=6200 $Y=1360
X8 10 M2_M1_CDNS_1 $T=7300 1510 0 90 $X=7170 $Y=1430
X9 9 M2_M1_CDNS_1 $T=7850 -2080 0 0 $X=7770 $Y=-2210
X10 10 M2_M1_CDNS_1 $T=9400 1510 0 90 $X=9270 $Y=1430
X11 6 M2_M1_CDNS_1 $T=9770 -2060 0 0 $X=9690 $Y=-2190
X12 1 M4_M3_CDNS_3 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X13 1 M4_M3_CDNS_3 $T=5110 3310 0 0 $X=5030 $Y=3060
X14 1 M3_M2_CDNS_6 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X15 1 M3_M2_CDNS_6 $T=5110 3310 0 0 $X=5030 $Y=3060
X16 11 M3_M2_CDNS_8 $T=1140 2170 0 90 $X=890 $Y=2090
X17 12 M3_M2_CDNS_8 $T=3910 970 0 0 $X=3830 $Y=720
X18 13 M3_M2_CDNS_8 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X19 11 M3_M2_CDNS_8 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X20 11 M3_M2_CDNS_8 $T=8100 2170 0 90 $X=7850 $Y=2090
X21 13 M3_M2_CDNS_8 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X22 12 M3_M2_CDNS_8 $T=9760 1890 0 0 $X=9680 $Y=1640
X23 11 M2_M1_CDNS_9 $T=1140 2170 0 90 $X=890 $Y=2090
X24 12 M2_M1_CDNS_9 $T=3910 970 0 0 $X=3830 $Y=720
X25 13 M2_M1_CDNS_9 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X26 11 M2_M1_CDNS_9 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X27 13 M2_M1_CDNS_9 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X28 12 M2_M1_CDNS_9 $T=9760 1890 0 0 $X=9680 $Y=1640
X29 1 M2_M1_CDNS_16 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X30 1 M2_M1_CDNS_16 $T=5110 3310 0 0 $X=5030 $Y=3060
X31 11 M2_M1_CDNS_16 $T=8100 2170 0 90 $X=7850 $Y=2090
X32 11 M1_PO_CDNS_17 $T=8100 2170 0 90 $X=7850 $Y=2070
X33 12 1 4 7 9 18 NAND2_1X_small $T=3680 -70 0 0 $X=3800 $Y=0
X34 3 1 4 7 INV_1X_small_layout $T=0 40 1 0 $X=0 $Y=-3760
X35 2 1 4 11 INV_1X_small_layout $T=0 0 0 0 $X=0 $Y=0
X36 6 1 4 8 INV_1X_small_layout $T=4800 40 1 0 $X=4800 $Y=-3760
X37 9 1 4 10 INV_1X_small_layout $T=6200 0 0 0 $X=6200 $Y=0
X38 13 1 4 6 INV_1X_small_layout $T=8600 40 1 0 $X=8600 $Y=-3760
X39 2 1 4 5 12 14 ph1p3_clk_part $T=1400 0 0 0 $X=1400 $Y=0
X40 2 1 4 8 13 15 ph1p3_clk_part $T=2400 40 1 0 $X=2400 $Y=-3760
X41 11 1 4 9 13 16 ph1p3_clk_part $T=6200 40 1 0 $X=6200 $Y=-3760
X42 11 1 4 10 12 17 ph1p3_clk_part $T=7600 0 0 0 $X=7600 $Y=0
X43 1 4 cellTmpl_CDNS_48 $T=1520 -100 1 0 $X=1400 $Y=-3760
.ends ph1p3_MSDFF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_49                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_49 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_49

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p1_MAC                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p1_MAC 40 38 37 32 42 43 33 39 34 35
+ 12 41 21 28 20 13 25 29 22 23
+ 30 17 26 27 36
** N=587 EP=25 FDC=1272
X0 1 M2_M1_CDNS_1 $T=13500 1730 0 90 $X=13370 $Y=1650
X1 2 M2_M1_CDNS_1 $T=26210 45120 0 0 $X=26130 $Y=44990
X2 3 M2_M1_CDNS_1 $T=27140 31160 0 0 $X=27060 $Y=31030
X3 4 M2_M1_CDNS_1 $T=27590 6180 0 0 $X=27510 $Y=6050
X4 5 M2_M1_CDNS_1 $T=27640 13250 0 0 $X=27560 $Y=13120
X5 6 M2_M1_CDNS_1 $T=27650 9990 0 0 $X=27570 $Y=9860
X6 7 M2_M1_CDNS_1 $T=27950 16370 0 90 $X=27820 $Y=16290
X7 8 M2_M1_CDNS_1 $T=35010 34430 0 0 $X=34930 $Y=34300
X8 9 M2_M1_CDNS_1 $T=35360 2150 0 90 $X=35230 $Y=2070
X9 10 M2_M1_CDNS_1 $T=36780 38020 0 0 $X=36700 $Y=37890
X10 4 M2_M1_CDNS_1 $T=40600 27670 0 0 $X=40520 $Y=27540
X11 11 M2_M1_CDNS_1 $T=42620 53320 0 0 $X=42540 $Y=53190
X12 12 M2_M1_CDNS_1 $T=46960 36680 0 0 $X=46880 $Y=36550
X13 13 M2_M1_CDNS_1 $T=47310 37030 0 0 $X=47230 $Y=36900
X14 14 M2_M1_CDNS_1 $T=50500 49780 0 90 $X=50370 $Y=49700
X15 15 M2_M1_CDNS_1 $T=50830 41480 0 270 $X=50700 $Y=41400
X16 5 M2_M1_CDNS_1 $T=50820 20570 0 0 $X=50740 $Y=20440
X17 16 M2_M1_CDNS_1 $T=50830 35140 0 0 $X=50750 $Y=35010
X18 7 M2_M1_CDNS_1 $T=50840 27900 0 0 $X=50760 $Y=27770
X19 3 M2_M1_CDNS_1 $T=50840 57040 0 0 $X=50760 $Y=56910
X20 17 M3_M2_CDNS_2 $T=13580 500 0 0 $X=13500 $Y=370
X21 1 M3_M2_CDNS_2 $T=21790 3100 0 0 $X=21710 $Y=2970
X22 17 M3_M2_CDNS_2 $T=23460 6480 0 0 $X=23380 $Y=6350
X23 18 M3_M2_CDNS_2 $T=25060 48910 0 0 $X=24980 $Y=48780
X24 10 M3_M2_CDNS_2 $T=27280 16600 0 0 $X=27200 $Y=16470
X25 19 M3_M2_CDNS_2 $T=27550 23950 0 0 $X=27470 $Y=23820
X26 3 M3_M2_CDNS_2 $T=31000 30620 0 90 $X=30870 $Y=30540
X27 18 M3_M2_CDNS_2 $T=31730 53970 0 0 $X=31650 $Y=53840
X28 8 M3_M2_CDNS_2 $T=36450 32450 0 0 $X=36370 $Y=32320
X29 8 M3_M2_CDNS_2 $T=37010 12970 0 0 $X=36930 $Y=12840
X30 4 M3_M2_CDNS_2 $T=37130 8320 0 90 $X=37000 $Y=8240
X31 4 M3_M2_CDNS_2 $T=37620 28370 0 0 $X=37540 $Y=28240
X32 13 M3_M2_CDNS_2 $T=39130 33810 0 0 $X=39050 $Y=33680
X33 14 M3_M2_CDNS_2 $T=39650 35610 0 90 $X=39520 $Y=35530
X34 16 M3_M2_CDNS_2 $T=41560 34270 0 0 $X=41480 $Y=34140
X35 20 M3_M2_CDNS_2 $T=45180 37600 0 0 $X=45100 $Y=37470
X36 21 M3_M2_CDNS_2 $T=47320 30390 0 0 $X=47240 $Y=30260
X37 21 M3_M2_CDNS_2 $T=47350 35870 0 0 $X=47270 $Y=35740
X38 5 M3_M2_CDNS_2 $T=47710 20800 0 0 $X=47630 $Y=20670
X39 7 M3_M2_CDNS_2 $T=47720 28200 0 0 $X=47640 $Y=28070
X40 12 M3_M2_CDNS_2 $T=47890 54000 0 0 $X=47810 $Y=53870
X41 22 M3_M2_CDNS_2 $T=47970 15770 0 0 $X=47890 $Y=15640
X42 3 M3_M2_CDNS_2 $T=49120 57660 0 90 $X=48990 $Y=57580
X43 23 M3_M2_CDNS_2 $T=50140 8430 0 0 $X=50060 $Y=8300
X44 24 M4_M3_CDNS_3 $T=14240 34180 0 0 $X=14160 $Y=33930
X45 2 M4_M3_CDNS_3 $T=14690 34260 0 0 $X=14610 $Y=34010
X46 16 M4_M3_CDNS_3 $T=27580 20920 0 0 $X=27500 $Y=20670
X47 11 M4_M3_CDNS_3 $T=29900 48890 0 0 $X=29820 $Y=48640
X48 19 M4_M3_CDNS_3 $T=30080 30230 0 90 $X=29830 $Y=30150
X49 10 M4_M3_CDNS_3 $T=30460 28380 0 90 $X=30210 $Y=28300
X50 10 M4_M3_CDNS_3 $T=30460 23030 0 0 $X=30380 $Y=22780
X51 19 M4_M3_CDNS_3 $T=30500 32130 0 0 $X=30420 $Y=31880
X52 5 M4_M3_CDNS_3 $T=33780 15450 0 0 $X=33700 $Y=15200
X53 7 M4_M3_CDNS_3 $T=35610 26220 0 0 $X=35530 $Y=25970
X54 19 M4_M3_CDNS_3 $T=36140 41490 0 0 $X=36060 $Y=41240
X55 13 M4_M3_CDNS_3 $T=37160 30260 0 0 $X=37080 $Y=30010
X56 25 M4_M3_CDNS_3 $T=37340 28940 0 0 $X=37260 $Y=28690
X57 19 M4_M3_CDNS_3 $T=38360 45240 0 0 $X=38280 $Y=44990
X58 9 M4_M3_CDNS_3 $T=40140 11980 0 0 $X=40060 $Y=11730
X59 9 M4_M3_CDNS_3 $T=40140 13750 0 0 $X=40060 $Y=13500
X60 6 M4_M3_CDNS_3 $T=41200 8070 0 0 $X=41120 $Y=7820
X61 26 M4_M3_CDNS_3 $T=42660 8560 0 0 $X=42580 $Y=8310
X62 12 M4_M3_CDNS_3 $T=45260 13780 0 0 $X=45180 $Y=13530
X63 12 M4_M3_CDNS_3 $T=46430 13570 0 0 $X=46350 $Y=13320
X64 12 M4_M3_CDNS_3 $T=46440 20680 0 0 $X=46360 $Y=20430
X65 12 M4_M3_CDNS_3 $T=46450 28020 0 0 $X=46370 $Y=27770
X66 27 M4_M3_CDNS_3 $T=48720 11410 0 0 $X=48640 $Y=11160
X67 27 M4_M3_CDNS_3 $T=48720 18740 0 0 $X=48640 $Y=18490
X68 27 M4_M3_CDNS_3 $T=48720 26060 0 0 $X=48640 $Y=25810
X69 27 M4_M3_CDNS_3 $T=48720 33370 0 0 $X=48640 $Y=33120
X70 27 M4_M3_CDNS_3 $T=48720 40760 0 0 $X=48640 $Y=40510
X71 27 M4_M3_CDNS_3 $T=48720 48010 0 0 $X=48640 $Y=47760
X72 27 M4_M3_CDNS_3 $T=48720 54650 0 0 $X=48640 $Y=54400
X73 15 M4_M3_CDNS_3 $T=50370 40700 0 90 $X=50120 $Y=40620
X74 14 M4_M3_CDNS_4 $T=31920 35650 0 90 $X=31670 $Y=35570
X75 8 M4_M3_CDNS_4 $T=32900 32450 0 90 $X=32650 $Y=32370
X76 20 M4_M3_CDNS_4 $T=33420 28560 0 0 $X=33340 $Y=28310
X77 28 M4_M3_CDNS_4 $T=33550 30080 0 0 $X=33470 $Y=29830
X78 25 M4_M3_CDNS_4 $T=33910 21000 0 0 $X=33830 $Y=20750
X79 29 M4_M3_CDNS_4 $T=35700 20190 0 0 $X=35620 $Y=19940
X80 22 M4_M3_CDNS_4 $T=36040 13890 0 0 $X=35960 $Y=13640
X81 3 M4_M3_CDNS_4 $T=36940 32400 0 0 $X=36860 $Y=32150
X82 5 M4_M3_CDNS_4 $T=37360 20060 0 0 $X=37280 $Y=19810
X83 22 M4_M3_CDNS_4 $T=40000 16980 0 90 $X=39750 $Y=16900
X84 5 M4_M3_CDNS_4 $T=40200 20060 0 90 $X=39950 $Y=19980
X85 23 M4_M3_CDNS_4 $T=40270 9670 0 90 $X=40020 $Y=9590
X86 7 M4_M3_CDNS_4 $T=40100 26260 0 0 $X=40020 $Y=26010
X87 3 M4_M3_CDNS_4 $T=42170 35070 0 90 $X=41920 $Y=34990
X88 12 M4_M3_CDNS_4 $T=47430 45810 0 0 $X=47350 $Y=45560
X89 24 M4_M3_CDNS_5 $T=13250 9080 0 0 $X=13170 $Y=8950
X90 24 M4_M3_CDNS_5 $T=13250 17420 0 0 $X=13170 $Y=17290
X91 24 M4_M3_CDNS_5 $T=13250 19900 0 0 $X=13170 $Y=19770
X92 2 M4_M3_CDNS_5 $T=13630 21000 0 0 $X=13550 $Y=20870
X93 18 M4_M3_CDNS_5 $T=24130 43430 0 0 $X=24050 $Y=43300
X94 11 M4_M3_CDNS_5 $T=27540 27470 0 0 $X=27460 $Y=27340
X95 18 M4_M3_CDNS_5 $T=27660 30880 0 0 $X=27580 $Y=30750
X96 17 M4_M3_CDNS_5 $T=29860 6490 0 0 $X=29780 $Y=6360
X97 30 M4_M3_CDNS_5 $T=30570 8500 0 90 $X=30440 $Y=8420
X98 23 M4_M3_CDNS_5 $T=33810 8340 0 0 $X=33730 $Y=8210
X99 13 M4_M3_CDNS_5 $T=34110 23130 0 0 $X=34030 $Y=23000
X100 30 M4_M3_CDNS_5 $T=34230 12140 0 0 $X=34150 $Y=12010
X101 15 M4_M3_CDNS_5 $T=35640 30080 0 0 $X=35560 $Y=29950
X102 20 M4_M3_CDNS_5 $T=36080 37590 0 90 $X=35950 $Y=37510
X103 5 M4_M3_CDNS_5 $T=36790 15500 0 0 $X=36710 $Y=15370
X104 16 M4_M3_CDNS_5 $T=36850 22810 0 0 $X=36770 $Y=22680
X105 4 M4_M3_CDNS_5 $T=37090 18980 0 0 $X=37010 $Y=18850
X106 4 M4_M3_CDNS_5 $T=37210 21640 0 0 $X=37130 $Y=21510
X107 1 M4_M3_CDNS_5 $T=37910 9490 0 0 $X=37830 $Y=9360
X108 1 M4_M3_CDNS_5 $T=40250 21000 0 0 $X=40170 $Y=20870
X109 26 M4_M3_CDNS_5 $T=40660 2660 0 0 $X=40580 $Y=2530
X110 12 M4_M3_CDNS_5 $T=46940 30240 0 0 $X=46860 $Y=30110
X111 21 M4_M3_CDNS_5 $T=47710 14100 0 0 $X=47630 $Y=13970
X112 21 M4_M3_CDNS_5 $T=47710 17150 0 0 $X=47630 $Y=17020
X113 6 M4_M3_CDNS_5 $T=50450 13720 0 180 $X=50370 $Y=13590
X114 24 M3_M2_CDNS_6 $T=14240 34180 0 0 $X=14160 $Y=33930
X115 14 M3_M2_CDNS_6 $T=27160 26930 0 0 $X=27080 $Y=26680
X116 16 M3_M2_CDNS_6 $T=27580 20920 0 0 $X=27500 $Y=20670
X117 8 M3_M2_CDNS_6 $T=32010 34020 0 90 $X=31760 $Y=33940
X118 30 M3_M2_CDNS_6 $T=33210 6090 0 90 $X=32960 $Y=6010
X119 28 M3_M2_CDNS_6 $T=34670 53910 0 0 $X=34590 $Y=53660
X120 13 M3_M2_CDNS_6 $T=37160 30260 0 0 $X=37080 $Y=30010
X121 17 M3_M2_CDNS_6 $T=37760 15780 0 0 $X=37680 $Y=15530
X122 30 M3_M2_CDNS_6 $T=37790 22530 0 0 $X=37710 $Y=22280
X123 29 M3_M2_CDNS_6 $T=37810 21110 0 0 $X=37730 $Y=20860
X124 19 M3_M2_CDNS_6 $T=38360 45240 0 0 $X=38280 $Y=44990
X125 9 M3_M2_CDNS_6 $T=40140 13750 0 0 $X=40060 $Y=13500
X126 1 M3_M2_CDNS_6 $T=40250 21000 0 0 $X=40170 $Y=20750
X127 12 M3_M2_CDNS_6 $T=46430 13570 0 0 $X=46350 $Y=13320
X128 12 M3_M2_CDNS_6 $T=46440 20680 0 0 $X=46360 $Y=20430
X129 12 M3_M2_CDNS_6 $T=46450 28020 0 0 $X=46370 $Y=27770
X130 27 M3_M2_CDNS_6 $T=48720 11410 0 0 $X=48640 $Y=11160
X131 27 M3_M2_CDNS_6 $T=48720 18740 0 0 $X=48640 $Y=18490
X132 27 M3_M2_CDNS_6 $T=48720 26060 0 0 $X=48640 $Y=25810
X133 27 M3_M2_CDNS_6 $T=48720 33370 0 0 $X=48640 $Y=33120
X134 27 M3_M2_CDNS_6 $T=48720 40760 0 0 $X=48640 $Y=40510
X135 27 M3_M2_CDNS_6 $T=48720 48010 0 0 $X=48640 $Y=47760
X136 27 M3_M2_CDNS_6 $T=48720 54650 0 0 $X=48640 $Y=54400
X137 12 M3_M2_CDNS_6 $T=49790 45580 0 90 $X=49540 $Y=45500
X138 6 M3_M2_CDNS_6 $T=50450 13720 0 180 $X=50370 $Y=13470
X139 2 M3_M2_CDNS_7 $T=14690 34260 0 0 $X=14610 $Y=34010
X140 11 M3_M2_CDNS_7 $T=29900 48890 0 0 $X=29820 $Y=48640
X141 19 M3_M2_CDNS_7 $T=30080 30230 0 90 $X=29830 $Y=30150
X142 10 M3_M2_CDNS_7 $T=30460 28380 0 90 $X=30210 $Y=28300
X143 10 M3_M2_CDNS_7 $T=30460 23030 0 0 $X=30380 $Y=22780
X144 19 M3_M2_CDNS_7 $T=30500 32130 0 0 $X=30420 $Y=31880
X145 5 M3_M2_CDNS_7 $T=33780 15450 0 0 $X=33700 $Y=15200
X146 7 M3_M2_CDNS_7 $T=35610 26220 0 0 $X=35530 $Y=25970
X147 19 M3_M2_CDNS_7 $T=36140 41490 0 0 $X=36060 $Y=41240
X148 25 M3_M2_CDNS_7 $T=37340 28940 0 0 $X=37260 $Y=28690
X149 9 M3_M2_CDNS_7 $T=40140 11980 0 0 $X=40060 $Y=11730
X150 6 M3_M2_CDNS_7 $T=41200 8070 0 0 $X=41120 $Y=7820
X151 26 M3_M2_CDNS_7 $T=42660 8560 0 0 $X=42580 $Y=8310
X152 12 M3_M2_CDNS_7 $T=45260 13780 0 0 $X=45180 $Y=13530
X153 12 M3_M2_CDNS_7 $T=46940 30240 0 0 $X=46860 $Y=29990
X154 15 M3_M2_CDNS_7 $T=50370 40700 0 90 $X=50120 $Y=40620
X155 31 M3_M2_CDNS_8 $T=22520 34180 0 0 $X=22440 $Y=33930
X156 15 M3_M2_CDNS_8 $T=27940 24310 0 0 $X=27860 $Y=24060
X157 18 M3_M2_CDNS_8 $T=31730 56230 0 0 $X=31650 $Y=55980
X158 21 M3_M2_CDNS_8 $T=39900 10160 0 90 $X=39650 $Y=10080
X159 21 M3_M2_CDNS_8 $T=39880 24880 0 0 $X=39800 $Y=24630
X160 21 M3_M2_CDNS_8 $T=39910 17530 0 0 $X=39830 $Y=17280
X161 13 M3_M2_CDNS_8 $T=45250 34520 0 0 $X=45170 $Y=34270
X162 21 M3_M2_CDNS_8 $T=47340 38170 0 90 $X=47090 $Y=38090
X163 21 M3_M2_CDNS_8 $T=47410 10180 0 0 $X=47330 $Y=9930
X164 21 M3_M2_CDNS_8 $T=47800 51890 0 90 $X=47550 $Y=51810
X165 21 M3_M2_CDNS_8 $T=47800 45070 0 0 $X=47720 $Y=44820
X166 21 M3_M2_CDNS_8 $T=48230 16850 0 0 $X=48150 $Y=16600
X167 21 M3_M2_CDNS_8 $T=48400 24170 0 0 $X=48320 $Y=23920
X168 24 M2_M1_CDNS_9 $T=14240 34180 0 0 $X=14160 $Y=33930
X169 31 M2_M1_CDNS_9 $T=22520 34180 0 0 $X=22440 $Y=33930
X170 15 M2_M1_CDNS_9 $T=27940 24310 0 0 $X=27860 $Y=24060
X171 18 M2_M1_CDNS_9 $T=31730 56230 0 0 $X=31650 $Y=55980
X172 19 M2_M1_CDNS_9 $T=38360 45240 0 0 $X=38280 $Y=44990
X173 13 M2_M1_CDNS_9 $T=45250 34520 0 0 $X=45170 $Y=34270
X174 14 M5_M4_CDNS_10 $T=27160 26930 0 0 $X=27080 $Y=26680
X175 14 M5_M4_CDNS_10 $T=31920 35650 0 90 $X=31670 $Y=35570
X176 8 M5_M4_CDNS_10 $T=32010 34020 0 90 $X=31760 $Y=33940
X177 8 M5_M4_CDNS_10 $T=32900 32450 0 90 $X=32650 $Y=32370
X178 30 M5_M4_CDNS_10 $T=33210 6090 0 90 $X=32960 $Y=6010
X179 20 M5_M4_CDNS_10 $T=33420 28560 0 0 $X=33340 $Y=28310
X180 28 M5_M4_CDNS_10 $T=33550 30080 0 0 $X=33470 $Y=29830
X181 25 M5_M4_CDNS_10 $T=33910 21000 0 0 $X=33830 $Y=20750
X182 28 M5_M4_CDNS_10 $T=34670 53910 0 0 $X=34590 $Y=53660
X183 29 M5_M4_CDNS_10 $T=35700 20190 0 0 $X=35620 $Y=19940
X184 22 M5_M4_CDNS_10 $T=36040 13890 0 0 $X=35960 $Y=13640
X185 3 M5_M4_CDNS_10 $T=36940 32400 0 0 $X=36860 $Y=32150
X186 5 M5_M4_CDNS_10 $T=37360 20060 0 0 $X=37280 $Y=19810
X187 17 M5_M4_CDNS_10 $T=37760 15780 0 0 $X=37680 $Y=15530
X188 30 M5_M4_CDNS_10 $T=37790 22530 0 0 $X=37710 $Y=22280
X189 29 M5_M4_CDNS_10 $T=37810 21110 0 0 $X=37730 $Y=20860
X190 22 M5_M4_CDNS_10 $T=40000 16980 0 90 $X=39750 $Y=16900
X191 5 M5_M4_CDNS_10 $T=40200 20060 0 90 $X=39950 $Y=19980
X192 23 M5_M4_CDNS_10 $T=40270 9670 0 90 $X=40020 $Y=9590
X193 7 M5_M4_CDNS_10 $T=40100 26260 0 0 $X=40020 $Y=26010
X194 3 M5_M4_CDNS_10 $T=42170 35070 0 90 $X=41920 $Y=34990
X195 12 M5_M4_CDNS_10 $T=47430 45810 0 0 $X=47350 $Y=45560
X196 12 M5_M4_CDNS_10 $T=49790 45580 0 90 $X=49540 $Y=45500
X197 14 M4_M3_CDNS_11 $T=27160 26930 0 0 $X=27080 $Y=26680
X198 8 M4_M3_CDNS_11 $T=32010 34020 0 90 $X=31760 $Y=33940
X199 30 M4_M3_CDNS_11 $T=33210 6090 0 90 $X=32960 $Y=6010
X200 28 M4_M3_CDNS_11 $T=34670 53910 0 0 $X=34590 $Y=53660
X201 17 M4_M3_CDNS_11 $T=37760 15780 0 0 $X=37680 $Y=15530
X202 30 M4_M3_CDNS_11 $T=37790 22530 0 0 $X=37710 $Y=22280
X203 29 M4_M3_CDNS_11 $T=37810 21110 0 0 $X=37730 $Y=20860
X204 12 M4_M3_CDNS_11 $T=49790 45580 0 90 $X=49540 $Y=45500
X205 30 M5_M4_CDNS_12 $T=30570 6460 0 0 $X=30490 $Y=6330
X206 28 M5_M4_CDNS_12 $T=32990 34750 0 0 $X=32910 $Y=34620
X207 28 M5_M4_CDNS_12 $T=34030 38880 0 0 $X=33950 $Y=38750
X208 28 M5_M4_CDNS_12 $T=34680 50390 0 0 $X=34600 $Y=50260
X209 25 M5_M4_CDNS_12 $T=34810 23910 0 0 $X=34730 $Y=23780
X210 28 M5_M4_CDNS_12 $T=35170 42160 0 0 $X=35090 $Y=42030
X211 30 M5_M4_CDNS_12 $T=35280 16530 0 0 $X=35200 $Y=16400
X212 20 M5_M4_CDNS_12 $T=36090 34240 0 0 $X=36010 $Y=34110
X213 15 M5_M4_CDNS_12 $T=36460 32950 0 0 $X=36380 $Y=32820
X214 17 M5_M4_CDNS_12 $T=37190 13870 0 0 $X=37110 $Y=13740
X215 23 M5_M4_CDNS_12 $T=37340 9680 0 0 $X=37260 $Y=9550
X216 26 M5_M4_CDNS_12 $T=37540 8130 0 0 $X=37460 $Y=8000
X217 1 M5_M4_CDNS_12 $T=38230 18800 0 90 $X=38100 $Y=18720
X218 7 M5_M4_CDNS_12 $T=38290 26230 0 90 $X=38160 $Y=26150
X219 1 M5_M4_CDNS_12 $T=39740 18800 0 90 $X=39610 $Y=18720
X220 26 M5_M4_CDNS_12 $T=39840 8560 0 90 $X=39710 $Y=8480
X221 6 M5_M4_CDNS_12 $T=47900 8080 0 0 $X=47820 $Y=7950
X222 6 M5_M4_CDNS_12 $T=49870 8100 0 0 $X=49790 $Y=7970
X223 15 M5_M4_CDNS_12 $T=49880 37370 0 0 $X=49800 $Y=37240
X224 21 M1_PO_CDNS_13 $T=47320 31410 0 0 $X=47220 $Y=31160
X225 12 M1_PO_CDNS_14 $T=47490 48870 0 0 $X=47390 $Y=48750
X226 21 M2_M1_CDNS_15 $T=47320 31410 0 0 $X=47240 $Y=31160
X227 14 M2_M1_CDNS_16 $T=27160 26930 0 0 $X=27080 $Y=26680
X228 16 M2_M1_CDNS_16 $T=27580 20920 0 0 $X=27500 $Y=20670
X229 30 M2_M1_CDNS_16 $T=33210 6090 0 90 $X=32960 $Y=6010
X230 13 M2_M1_CDNS_16 $T=37160 30260 0 0 $X=37080 $Y=30010
X231 21 M2_M1_CDNS_16 $T=39900 10160 0 90 $X=39650 $Y=10080
X232 21 M2_M1_CDNS_16 $T=39880 24880 0 0 $X=39800 $Y=24630
X233 21 M2_M1_CDNS_16 $T=39910 17530 0 0 $X=39830 $Y=17280
X234 9 M2_M1_CDNS_16 $T=40140 13750 0 0 $X=40060 $Y=13500
X235 1 M2_M1_CDNS_16 $T=40250 21000 0 0 $X=40170 $Y=20750
X236 12 M2_M1_CDNS_16 $T=46430 13570 0 0 $X=46350 $Y=13320
X237 12 M2_M1_CDNS_16 $T=46440 20680 0 0 $X=46360 $Y=20430
X238 12 M2_M1_CDNS_16 $T=46450 28020 0 0 $X=46370 $Y=27770
X239 21 M2_M1_CDNS_16 $T=47340 38170 0 90 $X=47090 $Y=38090
X240 21 M2_M1_CDNS_16 $T=47410 10180 0 0 $X=47330 $Y=9930
X241 21 M2_M1_CDNS_16 $T=47800 51890 0 90 $X=47550 $Y=51810
X242 21 M2_M1_CDNS_16 $T=47800 45070 0 0 $X=47720 $Y=44820
X243 21 M2_M1_CDNS_16 $T=48230 16850 0 0 $X=48150 $Y=16600
X244 21 M2_M1_CDNS_16 $T=48400 24170 0 0 $X=48320 $Y=23920
X245 27 M2_M1_CDNS_16 $T=48720 11410 0 0 $X=48640 $Y=11160
X246 27 M2_M1_CDNS_16 $T=48720 18740 0 0 $X=48640 $Y=18490
X247 27 M2_M1_CDNS_16 $T=48720 26060 0 0 $X=48640 $Y=25810
X248 27 M2_M1_CDNS_16 $T=48720 33370 0 0 $X=48640 $Y=33120
X249 27 M2_M1_CDNS_16 $T=48720 40760 0 0 $X=48640 $Y=40510
X250 27 M2_M1_CDNS_16 $T=48720 48010 0 0 $X=48640 $Y=47760
X251 27 M2_M1_CDNS_16 $T=48720 54650 0 0 $X=48640 $Y=54400
X252 6 M2_M1_CDNS_16 $T=50450 13720 0 180 $X=50370 $Y=13470
X253 30 M1_PO_CDNS_17 $T=33210 6090 0 90 $X=32960 $Y=5990
X254 21 M1_PO_CDNS_17 $T=39900 10160 0 90 $X=39650 $Y=10060
X255 21 M1_PO_CDNS_17 $T=39880 24880 0 0 $X=39780 $Y=24630
X256 21 M1_PO_CDNS_17 $T=39910 17530 0 0 $X=39810 $Y=17280
X257 12 M1_PO_CDNS_17 $T=46430 13570 0 0 $X=46330 $Y=13320
X258 12 M1_PO_CDNS_17 $T=46440 20680 0 0 $X=46340 $Y=20430
X259 12 M1_PO_CDNS_17 $T=46450 28020 0 0 $X=46350 $Y=27770
X260 21 M1_PO_CDNS_17 $T=47340 38170 0 90 $X=47090 $Y=38070
X261 21 M1_PO_CDNS_17 $T=47410 10180 0 0 $X=47310 $Y=9930
X262 21 M1_PO_CDNS_17 $T=47800 51890 0 90 $X=47550 $Y=51790
X263 21 M1_PO_CDNS_17 $T=47800 45070 0 0 $X=47700 $Y=44820
X264 21 M1_PO_CDNS_17 $T=48230 16850 0 0 $X=48130 $Y=16600
X265 21 M1_PO_CDNS_17 $T=48400 24170 0 0 $X=48300 $Y=23920
X266 32 27 33 34 35 36 37 38 39 24
+ 40 31 2 18 8 10 19 11 63 121
+ 110 127 50 148 131 93 147 149 62 59
+ 49 97 145 109 47 120 108 106 124 138
+ 81 84 144 82 91 45 55 119 80 92 multiplier $T=630 33200 0 0 $X=290 $Y=32980
X267 17 41 36 27 42 10 18 30 23 22
+ 25 13 20 28 11 19 2 29 8 24
+ 31 1 26 43 3 16 15 14 4 6
+ 5 7 9 44 171 170 175 174 163 173
+ 172 209 279 180 179 178 177 183 182 189
+ 188 187 186 165 164 167 166 169 168 10badder $T=-50850 53720 1 0 $X=-570 $Y=-60
X268 36 12 21 27 9 26 285 552 286 554
+ 288 284 289 282 283 287 290 ph1p3_MSDFF $T=37460 11020 0 0 $X=37460 $Y=7260
X269 36 12 21 27 1 17 294 555 295 557
+ 297 293 298 291 292 296 299 ph1p3_MSDFF $T=37460 18340 0 0 $X=37460 $Y=14580
X270 36 12 21 27 4 30 303 558 304 560
+ 306 302 307 300 301 305 308 ph1p3_MSDFF $T=37460 25660 0 0 $X=37460 $Y=21900
X271 36 12 21 27 6 23 312 561 313 563
+ 315 311 316 309 310 314 317 ph1p3_MSDFF $T=47700 11020 0 0 $X=47700 $Y=7260
X272 36 12 21 27 5 22 321 564 322 566
+ 324 320 325 318 319 323 326 ph1p3_MSDFF $T=47700 18340 0 0 $X=47700 $Y=14580
X273 36 12 21 27 7 29 330 567 331 569
+ 333 329 334 327 328 332 335 ph1p3_MSDFF $T=47700 25660 0 0 $X=47700 $Y=21900
X274 36 12 21 27 16 25 339 570 340 572
+ 342 338 343 336 337 341 344 ph1p3_MSDFF $T=47700 32980 0 0 $X=47700 $Y=29220
X275 36 12 21 27 15 13 348 573 349 575
+ 351 347 352 345 346 350 353 ph1p3_MSDFF $T=47700 40300 0 0 $X=47700 $Y=36540
X276 36 12 21 27 14 20 357 576 358 578
+ 360 356 361 354 355 359 362 ph1p3_MSDFF $T=47700 47620 0 0 $X=47700 $Y=43860
X277 36 12 21 27 3 28 366 579 367 581
+ 369 365 370 363 364 368 371 ph1p3_MSDFF $T=47700 54940 0 0 $X=47700 $Y=51180
X278 36 27 cellTmpl_CDNS_49 $T=47160 54840 1 0 $X=47040 $Y=51180
M0 285 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38240 $Y=8150 $dt=1
M1 288 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38240 $Y=13450 $dt=1
M2 294 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38240 $Y=15470 $dt=1
M3 297 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38240 $Y=20770 $dt=1
M4 303 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38240 $Y=22790 $dt=1
M5 306 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38240 $Y=28090 $dt=1
M6 282 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=39570 $Y=13480 $dt=1
M7 291 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=39570 $Y=20800 $dt=1
M8 300 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=39570 $Y=28120 $dt=1
M9 283 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=40570 $Y=8120 $dt=1
M10 292 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40570 $Y=15440 $dt=1
M11 301 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40570 $Y=22760 $dt=1
M12 284 12 9 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=40750 $Y=13480 $dt=1
M13 293 12 1 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=40750 $Y=20800 $dt=1
M14 302 12 4 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=40750 $Y=28120 $dt=1
M15 289 12 552 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=41750 $Y=8360 $dt=1
M16 298 12 555 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41750 $Y=15680 $dt=1
M17 307 12 558 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41750 $Y=23000 $dt=1
M18 286 284 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=41950 $Y=13390 $dt=1
M19 295 293 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=41950 $Y=20710 $dt=1
M20 304 302 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=41950 $Y=28030 $dt=1
M21 552 26 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=43040 $Y=8150 $dt=1
M22 555 17 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43040 $Y=15470 $dt=1
M23 558 30 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43040 $Y=22790 $dt=1
M24 286 285 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43190 $Y=13400 $dt=1
M25 295 294 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43190 $Y=20720 $dt=1
M26 304 303 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43190 $Y=28040 $dt=1
M27 287 288 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=44370 $Y=8120 $dt=1
M28 296 297 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44370 $Y=15440 $dt=1
M29 305 306 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44370 $Y=22760 $dt=1
M30 554 286 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44440 $Y=13450 $dt=1
M31 557 295 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44440 $Y=20770 $dt=1
M32 560 304 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=44440 $Y=28090 $dt=1
M33 289 288 286 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=45550 $Y=8360 $dt=1
M34 298 297 295 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=45550 $Y=15680 $dt=1
M35 307 306 304 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=45550 $Y=23000 $dt=1
M36 290 288 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=45770 $Y=13480 $dt=1
M37 299 297 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=45770 $Y=20800 $dt=1
M38 308 306 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=45770 $Y=28120 $dt=1
M39 26 289 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=46840 $Y=8150 $dt=1
M40 17 298 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=46840 $Y=15470 $dt=1
M41 30 307 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=46840 $Y=22790 $dt=1
M42 284 288 554 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46950 $Y=13480 $dt=1
M43 293 297 557 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46950 $Y=20800 $dt=1
M44 302 306 560 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=46950 $Y=28120 $dt=1
M45 312 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=48480 $Y=8150 $dt=1
M46 315 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48480 $Y=13450 $dt=1
M47 321 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48480 $Y=15470 $dt=1
M48 324 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48480 $Y=20770 $dt=1
M49 330 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48480 $Y=22790 $dt=1
M50 333 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48480 $Y=28090 $dt=1
M51 339 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48480 $Y=30110 $dt=1
M52 342 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48480 $Y=35410 $dt=1
M53 348 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48480 $Y=37430 $dt=1
M54 351 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48480 $Y=42730 $dt=1
M55 357 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48480 $Y=44750 $dt=1
M56 360 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48480 $Y=50050 $dt=1
M57 366 21 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48480 $Y=52070 $dt=1
M58 369 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48480 $Y=57370 $dt=1
M59 309 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=49810 $Y=13480 $dt=1
M60 318 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=49810 $Y=20800 $dt=1
M61 327 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=49810 $Y=28120 $dt=1
M62 336 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=49810 $Y=35440 $dt=1
M63 345 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=49810 $Y=42760 $dt=1
M64 354 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=49810 $Y=50080 $dt=1
M65 363 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=49810 $Y=57400 $dt=1
M66 310 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=50810 $Y=8120 $dt=1
M67 319 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50810 $Y=15440 $dt=1
M68 328 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50810 $Y=22760 $dt=1
M69 337 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50810 $Y=30080 $dt=1
M70 346 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50810 $Y=37400 $dt=1
M71 355 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50810 $Y=44720 $dt=1
M72 364 12 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50810 $Y=52040 $dt=1
M73 311 12 6 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=50990 $Y=13480 $dt=1
M74 320 12 5 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=50990 $Y=20800 $dt=1
M75 329 12 7 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=50990 $Y=28120 $dt=1
M76 338 12 16 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=50990 $Y=35440 $dt=1
M77 347 12 15 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=50990 $Y=42760 $dt=1
M78 356 12 14 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=50990 $Y=50080 $dt=1
M79 365 12 3 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=50990 $Y=57400 $dt=1
M80 316 12 561 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=51990 $Y=8360 $dt=1
M81 325 12 564 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51990 $Y=15680 $dt=1
M82 334 12 567 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51990 $Y=23000 $dt=1
M83 343 12 570 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51990 $Y=30320 $dt=1
M84 352 12 573 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51990 $Y=37640 $dt=1
M85 361 12 576 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51990 $Y=44960 $dt=1
M86 370 12 579 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51990 $Y=52280 $dt=1
M87 313 311 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52190 $Y=13390 $dt=1
M88 322 320 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52190 $Y=20710 $dt=1
M89 331 329 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52190 $Y=28030 $dt=1
M90 340 338 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52190 $Y=35350 $dt=1
M91 349 347 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52190 $Y=42670 $dt=1
M92 358 356 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52190 $Y=49990 $dt=1
M93 367 365 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=52190 $Y=57310 $dt=1
M94 561 23 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=53280 $Y=8150 $dt=1
M95 564 22 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53280 $Y=15470 $dt=1
M96 567 29 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53280 $Y=22790 $dt=1
M97 570 25 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53280 $Y=30110 $dt=1
M98 573 13 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53280 $Y=37430 $dt=1
M99 576 20 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53280 $Y=44750 $dt=1
M100 579 28 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53280 $Y=52070 $dt=1
M101 313 312 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53430 $Y=13400 $dt=1
M102 322 321 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53430 $Y=20720 $dt=1
M103 331 330 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53430 $Y=28040 $dt=1
M104 340 339 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53430 $Y=35360 $dt=1
M105 349 348 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53430 $Y=42680 $dt=1
M106 358 357 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53430 $Y=50000 $dt=1
M107 367 366 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=53430 $Y=57320 $dt=1
M108 314 315 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=54610 $Y=8120 $dt=1
M109 323 324 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=54610 $Y=15440 $dt=1
M110 332 333 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=54610 $Y=22760 $dt=1
M111 341 342 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=54610 $Y=30080 $dt=1
M112 350 351 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=54610 $Y=37400 $dt=1
M113 359 360 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=54610 $Y=44720 $dt=1
M114 368 369 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=54610 $Y=52040 $dt=1
M115 563 313 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=54680 $Y=13450 $dt=1
M116 566 322 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=54680 $Y=20770 $dt=1
M117 569 331 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=54680 $Y=28090 $dt=1
M118 572 340 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=54680 $Y=35410 $dt=1
M119 575 349 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=54680 $Y=42730 $dt=1
M120 578 358 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=54680 $Y=50050 $dt=1
M121 581 367 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=54680 $Y=57370 $dt=1
M122 316 315 313 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=55790 $Y=8360 $dt=1
M123 325 324 322 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=55790 $Y=15680 $dt=1
M124 334 333 331 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=55790 $Y=23000 $dt=1
M125 343 342 340 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=55790 $Y=30320 $dt=1
M126 352 351 349 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=55790 $Y=37640 $dt=1
M127 361 360 358 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=55790 $Y=44960 $dt=1
M128 370 369 367 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=55790 $Y=52280 $dt=1
M129 317 315 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56010 $Y=13480 $dt=1
M130 326 324 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56010 $Y=20800 $dt=1
M131 335 333 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56010 $Y=28120 $dt=1
M132 344 342 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56010 $Y=35440 $dt=1
M133 353 351 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56010 $Y=42760 $dt=1
M134 362 360 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56010 $Y=50080 $dt=1
M135 371 369 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=56010 $Y=57400 $dt=1
M136 23 316 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=57080 $Y=8150 $dt=1
M137 22 325 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=57080 $Y=15470 $dt=1
M138 29 334 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=57080 $Y=22790 $dt=1
M139 25 343 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=57080 $Y=30110 $dt=1
M140 13 352 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=57080 $Y=37430 $dt=1
M141 20 361 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=57080 $Y=44750 $dt=1
M142 28 370 36 36 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=57080 $Y=52070 $dt=1
M143 311 315 563 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57190 $Y=13480 $dt=1
M144 320 324 566 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57190 $Y=20800 $dt=1
M145 329 333 569 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57190 $Y=28120 $dt=1
M146 338 342 572 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57190 $Y=35440 $dt=1
M147 347 351 575 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57190 $Y=42760 $dt=1
M148 356 360 578 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57190 $Y=50080 $dt=1
M149 365 369 581 36 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=57190 $Y=57400 $dt=1
.ends ph2p1_MAC
