* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : MUX_4X                                       *
* Netlisted  : Thu Oct 24 16:36:29 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_3                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_3 S_source_0 D_drain_1 3 B
** N=5 EP=4 FDC=1
M0 D_drain_1 3 S_source_0 B g45p1svt L=4.5e-08 W=9.6e-07 AD=1.344e-13 AS=1.344e-13 PD=2.2e-06 PS=2.2e-06 fw=9.6e-07 sa=1.4e-07 sb=1.4e-07 sca=13.9449 scb=0.013907 scc=0.000385745 $X=0 $Y=0 $dt=1
.ends pmos1v_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_5                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_5 S_source_0 2 D_drain_1 4
** N=4 EP=4 FDC=1
M0 D_drain_1 2 S_source_0 4 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.72117 scb=0.00853087 scc=0.000206786 $X=0 $Y=0 $dt=0
.ends nmos1v_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_4X                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_4X A B Out S gnd! vdd!
** N=12 EP=6 FDC=12
X9 vdd! Out 7 vdd! pmos1v_CDNS_3 $T=5820 2540 0 270 $X=5620 $Y=2030
X15 gnd! S 4 gnd! nmos1v_CDNS_5 $T=750 890 0 0 $X=330 $Y=690
X16 gnd! 4 1 gnd! nmos1v_CDNS_5 $T=2140 890 0 0 $X=1720 $Y=690
X17 gnd! S 12 gnd! nmos1v_CDNS_5 $T=3070 890 0 0 $X=2650 $Y=690
X18 1 A 7 gnd! nmos1v_CDNS_5 $T=4000 890 0 0 $X=3580 $Y=690
X19 12 B 7 gnd! nmos1v_CDNS_5 $T=4930 890 0 0 $X=4510 $Y=690
X20 gnd! 7 Out gnd! nmos1v_CDNS_5 $T=6310 890 0 0 $X=5890 $Y=690
M0 4 S vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=17.2789 scb=0.0178533 scc=0.000435231 $X=750 $Y=2330 $dt=1
M1 2 4 vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=2140 $Y=2330 $dt=1
M2 11 S vdd! vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=3070 $Y=2330 $dt=1
M3 7 A 11 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=4000 $Y=2330 $dt=1
M4 7 B 2 vdd! g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7234 scb=0.0101098 scc=0.000278382 $X=4930 $Y=2330 $dt=1
.ends MUX_4X
