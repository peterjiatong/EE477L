* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : ph3_sytolic_array                            *
* Netlisted  : Sun Dec  8 17:46:28 2024                     *
* Pegasus Version: 22.21-s012 Fri Mar 10 17:36:33 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(g45n1svt) _nmos1v ndiff_conn(D) poly_conn(G) ndiff_conn(S) psubstrate(B)
*.DEVTMPLT 1 MP(g45p1svt) _pmos1v pdiff_conn(D) poly_conn(G) pdiff_conn(S) nwell_conn(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_1                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_1 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_2                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_2 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_3                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_3 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_4                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_4 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_4

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_5                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_5 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_5

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_6                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_6 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_6

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_7                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_7 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_7

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_8                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_8 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_8

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_9                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_9 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_9

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M5_M4_CDNS_10                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M5_M4_CDNS_10 1
** N=1 EP=1 FDC=0
.ends M5_M4_CDNS_10

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_11                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_11 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_11

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_12                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_12 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_12

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M4_M3_CDNS_13                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M4_M3_CDNS_13 1
** N=1 EP=1 FDC=0
.ends M4_M3_CDNS_13

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_14                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_14 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_14

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_15                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_15 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_15

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_16                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_16 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_16

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_17                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_17 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_17

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_18                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_18 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_18

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_new                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_new 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 3 M1_PO_CDNS_16 $T=1020 1750 0 90 $X=900 $Y=1650
X1 1 2 cellTmpl_CDNS_18 $T=50 150 0 0 $X=-70 $Y=10
M0 4 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.3086 scb=0.00950139 scc=0.000267597 $X=1140 $Y=930 $dt=0
.ends INV_1X_new

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_19                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_19 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_19

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_20                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_20 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_20

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_21                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_21 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_21

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND2_1X_small                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND2_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_16 $T=690 1680 0 90 $X=570 $Y=1580
X1 4 M1_PO_CDNS_16 $T=1930 1650 0 90 $X=1810 $Y=1550
X2 3 1 6 3 nmos1v_CDNS_19 $T=810 1000 0 0 $X=390 $Y=800
X3 6 4 5 3 nmos1v_CDNS_19 $T=2050 1000 0 0 $X=1630 $Y=800
X4 2 1 5 3 2 pmos1v_CDNS_20 $T=810 2440 0 0 $X=390 $Y=2240
X5 2 4 5 3 2 pmos1v_CDNS_20 $T=2050 2450 0 0 $X=1630 $Y=2250
X6 2 3 cellTmpl_CDNS_21 $T=240 210 0 0 $X=120 $Y=70
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=810 $Y=1000 $dt=0
M1 5 4 6 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=10.5213 scb=0.00984539 scc=0.000291491 $X=2050 $Y=1000 $dt=0
.ends NAND2_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: AND                                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt AND 1 2 3 4 5 6
*.DEVICECLIMB
** N=7 EP=6 FDC=3
X0 2 3 6 5 INV_1X_new $T=2480 -10 0 0 $X=2410 $Y=0
X1 1 2 3 4 6 7 NAND2_1X_small $T=-110 -70 0 0 $X=10 $Y=0
.ends AND

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_22                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_22 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_22

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1_PO_CDNS_23                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1_PO_CDNS_23 1
** N=1 EP=1 FDC=0
.ends M1_PO_CDNS_23

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M3_M2_CDNS_24                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M3_M2_CDNS_24 1
** N=1 EP=1 FDC=0
.ends M3_M2_CDNS_24

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_25                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_25 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_25

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M2_M1_CDNS_26                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M2_M1_CDNS_26 1
** N=1 EP=1 FDC=0
.ends M2_M1_CDNS_26

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_27                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_27 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_27

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_28                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_28 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_28

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_29                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_29 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_29

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR_small                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR_small 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=9
X0 1 M2_M1_CDNS_8 $T=350 1340 0 90 $X=220 $Y=1260
X1 6 M2_M1_CDNS_8 $T=5510 3180 0 90 $X=5380 $Y=3100
X2 6 M2_M1_CDNS_8 $T=6740 3180 0 90 $X=6610 $Y=3100
X3 1 M1_PO_CDNS_16 $T=580 1660 0 90 $X=460 $Y=1560
X4 4 M1_PO_CDNS_16 $T=1990 1480 0 90 $X=1870 $Y=1380
X5 4 M1_PO_CDNS_22 $T=5990 1680 0 90 $X=5790 $Y=1580
X6 1 M1_PO_CDNS_22 $T=7100 1350 0 90 $X=6900 $Y=1250
X7 7 M1_PO_CDNS_23 $T=3070 1660 0 90 $X=2870 $Y=1560
X8 8 M1_PO_CDNS_23 $T=4410 1540 0 90 $X=4210 $Y=1440
X9 8 M3_M2_CDNS_24 $T=1210 1540 0 90 $X=1010 $Y=1440
X10 8 M3_M2_CDNS_24 $T=4410 1540 0 90 $X=4210 $Y=1440
X11 8 M2_M1_CDNS_25 $T=1210 1540 0 90 $X=1010 $Y=1440
X12 4 M2_M1_CDNS_25 $T=1820 1880 0 90 $X=1620 $Y=1780
X13 8 M2_M1_CDNS_25 $T=4410 1540 0 90 $X=4210 $Y=1440
X14 4 M2_M1_CDNS_26 $T=5990 1680 0 90 $X=5790 $Y=1580
X15 1 M2_M1_CDNS_26 $T=7100 1350 0 90 $X=6900 $Y=1250
X16 2 3 cellTmpl_CDNS_27 $T=120 140 0 0 $X=0 $Y=0
X17 2 1 8 3 2 pmos1v_CDNS_28 $T=700 2180 0 0 $X=280 $Y=1980
X18 2 4 7 3 2 pmos1v_CDNS_28 $T=2110 2170 0 0 $X=1690 $Y=1970
X19 2 7 6 3 2 pmos1v_CDNS_28 $T=3270 2160 0 0 $X=2850 $Y=1960
X20 2 8 6 3 2 pmos1v_CDNS_28 $T=4610 2160 0 0 $X=4190 $Y=1960
X21 6 4 5 3 2 pmos1v_CDNS_28 $T=6140 2120 0 0 $X=5720 $Y=1920
X22 6 1 5 3 2 pmos1v_CDNS_28 $T=7250 2160 0 0 $X=6830 $Y=1960
X23 3 1 8 3 nmos1v_CDNS_29 $T=700 590 0 0 $X=280 $Y=390
X24 3 4 7 3 nmos1v_CDNS_29 $T=2110 580 0 0 $X=1690 $Y=380
X25 3 7 9 3 nmos1v_CDNS_29 $T=3270 580 0 0 $X=2850 $Y=380
X26 9 8 5 3 nmos1v_CDNS_29 $T=4610 580 0 0 $X=4190 $Y=380
X27 3 4 10 3 nmos1v_CDNS_29 $T=6140 600 0 0 $X=5720 $Y=400
X28 10 1 5 3 nmos1v_CDNS_29 $T=7250 650 0 0 $X=6830 $Y=450
M0 8 1 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.45462 scb=0.00478425 scc=6.8709e-05 $X=700 $Y=590 $dt=0
M1 7 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=2110 $Y=580 $dt=0
M2 9 7 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=3270 $Y=580 $dt=0
M3 5 8 9 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.34996 scb=0.00460723 scc=6.29421e-05 $X=4610 $Y=580 $dt=0
M4 10 4 3 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.56294 scb=0.00496757 scc=7.49928e-05 $X=6140 $Y=600 $dt=0
M5 5 1 10 3 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=7250 $Y=650 $dt=0
M6 7 4 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.1869 scb=0.0086398 scc=0.00051649 $X=2110 $Y=2170 $dt=1
M7 6 7 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3270 $Y=2160 $dt=1
M8 6 8 2 2 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4610 $Y=2160 $dt=1
.ends XOR_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: half_adder                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt half_adder 1 2 3 4 5 6 8 9 13
*.DEVICECLIMB
** N=13 EP=9 FDC=12
X0 4 M3_M2_CDNS_1 $T=6750 2480 0 0 $X=6670 $Y=2230
X1 4 M3_M2_CDNS_1 $T=9120 2880 0 0 $X=9040 $Y=2630
X2 4 M2_M1_CDNS_9 $T=6750 2480 0 0 $X=6670 $Y=2230
X3 4 M2_M1_CDNS_9 $T=9120 2880 0 0 $X=9040 $Y=2630
X4 4 M1_PO_CDNS_14 $T=6750 2480 0 0 $X=6650 $Y=2230
X5 4 M1_PO_CDNS_14 $T=9120 2880 0 0 $X=9020 $Y=2630
X6 1 3 2 4 6 9 AND $T=7790 0 0 0 $X=7800 $Y=0
X7 1 3 2 4 5 13 7 8 10 11 XOR_small $T=0 0 0 0 $X=0 $Y=0
.ends half_adder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_33                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_33 1 2
*.DEVICECLIMB
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_33

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_1X_small                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_1X_small 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=-310 120 0 0 $X=-430 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1000 $Y=830 $dt=0
M1 4 5 6 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=12.2783 scb=0.012115 scc=0.000626647 $X=1210 $Y=830 $dt=0
.ends NAND_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: NAND_2X_small1                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt NAND_2X_small1 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 2 cellTmpl_CDNS_33 $T=130 160 0 0 $X=10 $Y=20
M0 6 4 2 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=7.66878 scb=0.00580736 scc=7.77234e-05 $X=940 $Y=890 $dt=0
M1 3 5 6 2 g45n1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=11.676 scb=0.0124835 scc=0.000479408 $X=940 $Y=1100 $dt=0
.ends NAND_2X_small1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_39                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_39 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_39

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: XOR1                                            *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt XOR1 1 2 3 4 5 6 7 8 9 10
*.DEVICECLIMB
** N=10 EP=10 FDC=6
X0 6 M2_M1_CDNS_8 $T=1210 1480 0 90 $X=1080 $Y=1400
X1 7 M2_M1_CDNS_8 $T=2250 1860 0 90 $X=2120 $Y=1780
X2 6 M2_M1_CDNS_8 $T=2950 1480 0 90 $X=2820 $Y=1400
X3 8 M2_M1_CDNS_8 $T=3370 650 0 0 $X=3290 $Y=520
X4 9 M2_M1_CDNS_8 $T=3370 3080 0 0 $X=3290 $Y=2950
X5 9 M2_M1_CDNS_8 $T=3930 3080 0 0 $X=3850 $Y=2950
X6 7 M2_M1_CDNS_8 $T=4680 1860 0 90 $X=4550 $Y=1780
X7 9 M2_M1_CDNS_8 $T=4890 3070 0 0 $X=4810 $Y=2940
X8 8 M2_M1_CDNS_8 $T=5840 640 0 0 $X=5760 $Y=510
X9 9 M2_M1_CDNS_8 $T=6260 3080 0 0 $X=6180 $Y=2950
X10 6 M1_PO_CDNS_16 $T=4020 1500 0 90 $X=3900 $Y=1400
X11 7 M1_PO_CDNS_16 $T=5020 1730 0 90 $X=4900 $Y=1630
X12 2 3 6 2 nmos1v_CDNS_19 $T=830 840 0 0 $X=410 $Y=640
X13 2 4 7 2 nmos1v_CDNS_19 $T=1790 840 0 0 $X=1370 $Y=640
X14 1 3 6 2 1 pmos1v_CDNS_20 $T=830 2320 0 0 $X=410 $Y=2120
X15 1 4 7 2 1 pmos1v_CDNS_20 $T=1790 2320 0 0 $X=1370 $Y=2120
X16 1 4 9 2 1 pmos1v_CDNS_28 $T=3120 2080 0 0 $X=2700 $Y=1880
X17 9 6 5 2 1 pmos1v_CDNS_28 $T=4090 2140 0 0 $X=3670 $Y=1940
X18 9 7 5 2 1 pmos1v_CDNS_28 $T=5050 2140 0 0 $X=4630 $Y=1940
X19 1 3 9 2 1 pmos1v_CDNS_28 $T=6010 2140 0 0 $X=5590 $Y=1940
X20 2 4 8 2 nmos1v_CDNS_29 $T=3120 780 0 0 $X=2700 $Y=580
X21 10 6 5 2 nmos1v_CDNS_29 $T=4090 760 0 0 $X=3670 $Y=560
X22 10 7 2 2 nmos1v_CDNS_29 $T=5050 770 0 0 $X=4630 $Y=570
X23 8 3 5 2 nmos1v_CDNS_29 $T=6010 770 0 0 $X=5590 $Y=570
X24 1 2 cellTmpl_CDNS_39 $T=180 120 0 0 $X=60 $Y=-20
M0 6 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=830 $Y=840 $dt=0
M1 7 4 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1790 $Y=840 $dt=0
M2 8 4 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=3120 $Y=780 $dt=0
M3 5 6 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4126 scb=0.0095497 scc=0.000351079 $X=4090 $Y=760 $dt=0
M4 2 7 10 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=5050 $Y=770 $dt=0
M5 5 3 8 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=6010 $Y=770 $dt=0
.ends XOR1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: full_adder1_small                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt full_adder1_small 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 22 23
*.DEVICECLIMB
** N=23 EP=16 FDC=18
X0 1 M3_M2_CDNS_1 $T=590 2080 0 90 $X=340 $Y=2000
X1 3 M3_M2_CDNS_1 $T=2300 3150 0 90 $X=2050 $Y=3070
X2 1 M3_M2_CDNS_1 $T=17380 1890 0 0 $X=17300 $Y=1640
X3 3 M3_M2_CDNS_1 $T=19040 3010 0 0 $X=18960 $Y=2760
X4 8 M3_M2_CDNS_4 $T=6970 950 0 0 $X=6890 $Y=820
X5 8 M3_M2_CDNS_4 $T=14100 570 0 90 $X=13970 $Y=490
X6 8 M2_M1_CDNS_8 $T=6580 1900 0 0 $X=6500 $Y=1770
X7 9 M2_M1_CDNS_8 $T=15190 1730 0 90 $X=15060 $Y=1650
X8 1 M2_M1_CDNS_9 $T=590 2080 0 90 $X=340 $Y=2000
X9 3 M2_M1_CDNS_9 $T=2300 3150 0 90 $X=2050 $Y=3070
X10 1 M2_M1_CDNS_9 $T=17380 1890 0 0 $X=17300 $Y=1640
X11 3 M2_M1_CDNS_9 $T=19040 3010 0 0 $X=18960 $Y=2760
X12 1 M1_PO_CDNS_14 $T=590 2080 0 90 $X=340 $Y=1980
X13 3 M1_PO_CDNS_14 $T=2300 3150 0 90 $X=2050 $Y=3050
X14 1 M1_PO_CDNS_14 $T=17380 1890 0 0 $X=17280 $Y=1640
X15 3 M1_PO_CDNS_14 $T=19040 3010 0 0 $X=18940 $Y=2760
X16 8 M1_PO_CDNS_15 $T=8510 1970 0 0 $X=8410 $Y=1720
X17 8 M1_PO_CDNS_15 $T=16110 1570 0 0 $X=16010 $Y=1320
X18 9 M1_PO_CDNS_15 $T=20260 1840 0 0 $X=20160 $Y=1590
X19 1 M1_PO_CDNS_16 $T=690 1610 0 0 $X=590 $Y=1490
X20 3 M1_PO_CDNS_16 $T=1650 1990 0 0 $X=1550 $Y=1870
X21 5 M1_PO_CDNS_16 $T=7590 1960 0 0 $X=7490 $Y=1840
X22 10 M1_PO_CDNS_16 $T=19320 1680 0 0 $X=19220 $Y=1560
X23 8 M2_M1_CDNS_17 $T=8510 1970 0 0 $X=8430 $Y=1720
X24 8 M2_M1_CDNS_17 $T=16110 1570 0 0 $X=16030 $Y=1320
X25 9 M2_M1_CDNS_17 $T=20260 1840 0 0 $X=20180 $Y=1590
X26 2 4 1 10 3 20 NAND_1X_small $T=16970 30 0 0 $X=16540 $Y=10
X27 2 4 9 7 10 21 NAND_1X_small $T=19810 30 0 0 $X=19380 $Y=10
X28 2 4 9 5 8 19 NAND_2X_small1 $T=13690 -10 0 0 $X=13700 $Y=10
X29 2 4 1 3 8 11 12 15 22 16 XOR1 $T=-40 30 0 0 $X=20 $Y=10
X30 2 4 5 8 6 13 14 17 23 18 XOR1 $T=6800 30 0 0 $X=6860 $Y=10
.ends full_adder1_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: multiplier                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt multiplier 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
** N=238 EP=50 FDC=456
X0 2 M3_M2_CDNS_1 $T=160 15480 0 0 $X=80 $Y=15230
X1 2 M3_M2_CDNS_1 $T=160 21130 0 0 $X=80 $Y=20880
X2 2 M3_M2_CDNS_1 $T=170 9270 0 0 $X=90 $Y=9020
X3 2 M3_M2_CDNS_1 $T=170 13790 0 0 $X=90 $Y=13540
X4 19 M3_M2_CDNS_1 $T=500 8210 0 0 $X=420 $Y=7960
X5 1 M3_M2_CDNS_1 $T=1350 15570 0 0 $X=1270 $Y=15320
X6 1 M3_M2_CDNS_1 $T=1360 13320 0 0 $X=1280 $Y=13070
X7 20 M3_M2_CDNS_1 $T=4380 23070 0 90 $X=4130 $Y=22990
X8 21 M3_M2_CDNS_1 $T=4340 15320 0 0 $X=4260 $Y=15070
X9 22 M3_M2_CDNS_1 $T=5400 21130 0 0 $X=5320 $Y=20880
X10 7 M3_M2_CDNS_1 $T=5740 15570 0 0 $X=5660 $Y=15320
X11 7 M3_M2_CDNS_1 $T=5750 13320 0 0 $X=5670 $Y=13070
X12 19 M3_M2_CDNS_1 $T=6590 5910 0 0 $X=6510 $Y=5660
X13 23 M3_M2_CDNS_1 $T=7520 22860 0 0 $X=7440 $Y=22610
X14 23 M3_M2_CDNS_1 $T=7960 21030 0 0 $X=7880 $Y=20780
X15 24 M3_M2_CDNS_1 $T=8730 15340 0 0 $X=8650 $Y=15090
X16 8 M3_M2_CDNS_1 $T=8980 17010 0 0 $X=8900 $Y=16760
X17 8 M3_M2_CDNS_1 $T=10140 15570 0 0 $X=10060 $Y=15320
X18 8 M3_M2_CDNS_1 $T=10150 13320 0 0 $X=10070 $Y=13070
X19 25 M3_M2_CDNS_1 $T=12100 19160 0 0 $X=12020 $Y=18910
X20 20 M3_M2_CDNS_1 $T=12260 20780 0 0 $X=12180 $Y=20530
X21 26 M3_M2_CDNS_1 $T=13150 15340 0 0 $X=13070 $Y=15090
X22 27 M3_M2_CDNS_1 $T=14690 20780 0 0 $X=14610 $Y=20530
X23 28 M3_M2_CDNS_1 $T=15670 8330 0 0 $X=15590 $Y=8080
X24 29 M3_M2_CDNS_1 $T=16600 750 0 0 $X=16520 $Y=500
X25 27 M3_M2_CDNS_1 $T=17570 22850 0 0 $X=17490 $Y=22600
X26 30 M3_M2_CDNS_1 $T=22230 22840 0 0 $X=22150 $Y=22590
X27 30 M3_M2_CDNS_1 $T=28820 20830 0 0 $X=28740 $Y=20580
X28 31 M3_M2_CDNS_1 $T=35370 22940 0 0 $X=35290 $Y=22690
X29 2 M2_M1_CDNS_2 $T=160 15480 0 0 $X=80 $Y=15230
X30 2 M2_M1_CDNS_2 $T=160 21130 0 0 $X=80 $Y=20880
X31 2 M2_M1_CDNS_2 $T=170 9270 0 0 $X=90 $Y=9020
X32 2 M2_M1_CDNS_2 $T=170 13790 0 0 $X=90 $Y=13540
X33 19 M2_M1_CDNS_2 $T=500 8210 0 0 $X=420 $Y=7960
X34 20 M2_M1_CDNS_2 $T=4380 23070 0 90 $X=4130 $Y=22990
X35 21 M2_M1_CDNS_2 $T=4340 15320 0 0 $X=4260 $Y=15070
X36 22 M2_M1_CDNS_2 $T=5400 21130 0 0 $X=5320 $Y=20880
X37 24 M2_M1_CDNS_2 $T=8730 15340 0 0 $X=8650 $Y=15090
X38 25 M2_M1_CDNS_2 $T=12100 19160 0 0 $X=12020 $Y=18910
X39 26 M2_M1_CDNS_2 $T=13150 15340 0 0 $X=13070 $Y=15090
X40 27 M2_M1_CDNS_2 $T=17570 22850 0 0 $X=17490 $Y=22600
X41 30 M2_M1_CDNS_2 $T=22230 22840 0 0 $X=22150 $Y=22590
X42 30 M2_M1_CDNS_2 $T=28820 20830 0 0 $X=28740 $Y=20580
X43 31 M2_M1_CDNS_2 $T=35370 22940 0 0 $X=35290 $Y=22690
X44 32 M2_M1_CDNS_2 $T=46340 18970 0 0 $X=46260 $Y=18720
X45 33 M4_M3_CDNS_3 $T=34850 16990 0 0 $X=34770 $Y=16740
X46 21 M3_M2_CDNS_4 $T=4340 13390 0 0 $X=4260 $Y=13260
X47 22 M3_M2_CDNS_4 $T=7370 12440 0 0 $X=7290 $Y=12310
X48 22 M3_M2_CDNS_4 $T=8600 9080 0 0 $X=8520 $Y=8950
X49 8 M3_M2_CDNS_4 $T=10370 18740 0 0 $X=10290 $Y=18610
X50 25 M3_M2_CDNS_4 $T=13190 12020 0 0 $X=13110 $Y=11890
X51 34 M3_M2_CDNS_4 $T=19690 2880 0 90 $X=19560 $Y=2800
X52 35 M3_M2_CDNS_4 $T=26840 17540 0 90 $X=26710 $Y=17460
X53 31 M3_M2_CDNS_4 $T=35760 21100 0 0 $X=35680 $Y=20970
X54 30 M5_M4_CDNS_5 $T=34220 19150 0 0 $X=34140 $Y=18900
X55 33 M5_M4_CDNS_5 $T=34850 16990 0 0 $X=34770 $Y=16740
X56 30 M4_M3_CDNS_6 $T=28820 19250 0 0 $X=28740 $Y=19000
X57 30 M4_M3_CDNS_6 $T=34220 19150 0 0 $X=34140 $Y=18900
X58 1 M3_M2_CDNS_7 $T=1390 21140 0 0 $X=1310 $Y=20890
X59 7 M3_M2_CDNS_7 $T=4510 16920 0 0 $X=4430 $Y=16670
X60 36 M3_M2_CDNS_7 $T=8750 8160 0 0 $X=8670 $Y=7910
X61 37 M3_M2_CDNS_7 $T=10750 19470 0 0 $X=10670 $Y=19220
X62 38 M3_M2_CDNS_7 $T=11680 11800 0 0 $X=11600 $Y=11550
X63 35 M3_M2_CDNS_7 $T=13170 22790 0 0 $X=13090 $Y=22540
X64 11 M3_M2_CDNS_7 $T=13290 16990 0 0 $X=13210 $Y=16740
X65 11 M3_M2_CDNS_7 $T=14530 13310 0 0 $X=14450 $Y=13060
X66 11 M3_M2_CDNS_7 $T=14530 15600 0 0 $X=14450 $Y=15350
X67 38 M3_M2_CDNS_7 $T=22150 6400 0 0 $X=22070 $Y=6150
X68 39 M3_M2_CDNS_7 $T=24490 750 0 0 $X=24410 $Y=500
X69 40 M3_M2_CDNS_7 $T=26370 19410 0 0 $X=26290 $Y=19160
X70 33 M3_M2_CDNS_7 $T=26600 23000 0 0 $X=26520 $Y=22750
X71 30 M3_M2_CDNS_7 $T=28820 19250 0 0 $X=28740 $Y=19000
X72 41 M3_M2_CDNS_7 $T=29280 19170 0 0 $X=29200 $Y=18920
X73 37 M3_M2_CDNS_7 $T=33860 19960 0 90 $X=33610 $Y=19880
X74 30 M3_M2_CDNS_7 $T=34220 19150 0 0 $X=34140 $Y=18900
X75 42 M3_M2_CDNS_7 $T=35970 2380 0 0 $X=35890 $Y=2130
X76 41 M3_M2_CDNS_7 $T=39640 17490 0 0 $X=39560 $Y=17240
X77 28 M3_M2_CDNS_7 $T=43850 8260 0 0 $X=43770 $Y=8010
X78 29 M3_M2_CDNS_7 $T=43880 660 0 0 $X=43800 $Y=410
X79 32 M3_M2_CDNS_7 $T=46340 18970 0 0 $X=46260 $Y=18720
X80 2 M2_M1_CDNS_8 $T=170 4730 0 0 $X=90 $Y=4600
X81 2 M2_M1_CDNS_8 $T=180 890 0 0 $X=100 $Y=760
X82 43 M2_M1_CDNS_8 $T=4340 11800 0 0 $X=4260 $Y=11670
X83 39 M2_M1_CDNS_8 $T=8880 12210 0 0 $X=8800 $Y=12080
X84 44 M2_M1_CDNS_8 $T=13420 4530 0 0 $X=13340 $Y=4400
X85 45 M2_M1_CDNS_8 $T=17560 15460 0 0 $X=17480 $Y=15330
X86 34 M2_M1_CDNS_8 $T=21930 4780 0 0 $X=21850 $Y=4650
X87 46 M2_M1_CDNS_8 $T=29730 11900 0 0 $X=29650 $Y=11770
X88 47 M2_M1_CDNS_8 $T=31310 15530 0 0 $X=31230 $Y=15400
X89 48 M2_M1_CDNS_8 $T=35410 9580 0 0 $X=35330 $Y=9450
X90 49 M2_M1_CDNS_8 $T=41980 11840 0 0 $X=41900 $Y=11710
X91 42 M2_M1_CDNS_8 $T=43890 4790 0 0 $X=43810 $Y=4660
X92 1 M2_M1_CDNS_9 $T=1350 15570 0 0 $X=1270 $Y=15320
X93 1 M2_M1_CDNS_9 $T=1360 13320 0 0 $X=1280 $Y=13070
X94 1 M2_M1_CDNS_9 $T=1390 21140 0 0 $X=1310 $Y=20890
X95 7 M2_M1_CDNS_9 $T=4510 16920 0 0 $X=4430 $Y=16670
X96 7 M2_M1_CDNS_9 $T=5740 15570 0 0 $X=5660 $Y=15320
X97 7 M2_M1_CDNS_9 $T=5750 13320 0 0 $X=5670 $Y=13070
X98 19 M2_M1_CDNS_9 $T=6590 5910 0 0 $X=6510 $Y=5660
X99 23 M2_M1_CDNS_9 $T=7520 22860 0 0 $X=7440 $Y=22610
X100 23 M2_M1_CDNS_9 $T=7960 21030 0 0 $X=7880 $Y=20780
X101 36 M2_M1_CDNS_9 $T=8750 8160 0 0 $X=8670 $Y=7910
X102 8 M2_M1_CDNS_9 $T=8980 17010 0 0 $X=8900 $Y=16760
X103 8 M2_M1_CDNS_9 $T=10140 15570 0 0 $X=10060 $Y=15320
X104 8 M2_M1_CDNS_9 $T=10150 13320 0 0 $X=10070 $Y=13070
X105 8 M2_M1_CDNS_9 $T=10370 18740 0 0 $X=10290 $Y=18490
X106 37 M2_M1_CDNS_9 $T=10750 19470 0 0 $X=10670 $Y=19220
X107 38 M2_M1_CDNS_9 $T=11680 11800 0 0 $X=11600 $Y=11550
X108 20 M2_M1_CDNS_9 $T=12260 20780 0 0 $X=12180 $Y=20530
X109 35 M2_M1_CDNS_9 $T=13170 22790 0 0 $X=13090 $Y=22540
X110 11 M2_M1_CDNS_9 $T=13290 16990 0 0 $X=13210 $Y=16740
X111 11 M2_M1_CDNS_9 $T=14530 13310 0 0 $X=14450 $Y=13060
X112 11 M2_M1_CDNS_9 $T=14530 15600 0 0 $X=14450 $Y=15350
X113 27 M2_M1_CDNS_9 $T=14690 20780 0 0 $X=14610 $Y=20530
X114 28 M2_M1_CDNS_9 $T=15670 8330 0 0 $X=15590 $Y=8080
X115 29 M2_M1_CDNS_9 $T=16600 750 0 0 $X=16520 $Y=500
X116 38 M2_M1_CDNS_9 $T=22150 6400 0 0 $X=22070 $Y=6150
X117 39 M2_M1_CDNS_9 $T=24490 750 0 0 $X=24410 $Y=500
X118 40 M2_M1_CDNS_9 $T=26370 19410 0 0 $X=26290 $Y=19160
X119 33 M2_M1_CDNS_9 $T=26600 23000 0 0 $X=26520 $Y=22750
X120 30 M2_M1_CDNS_9 $T=28820 19250 0 0 $X=28740 $Y=19000
X121 41 M2_M1_CDNS_9 $T=29280 19170 0 0 $X=29200 $Y=18920
X122 37 M2_M1_CDNS_9 $T=33860 19960 0 90 $X=33610 $Y=19880
X123 30 M2_M1_CDNS_9 $T=34220 19150 0 0 $X=34140 $Y=18900
X124 31 M2_M1_CDNS_9 $T=35760 21100 0 0 $X=35680 $Y=20850
X125 42 M2_M1_CDNS_9 $T=35970 2380 0 0 $X=35890 $Y=2130
X126 41 M2_M1_CDNS_9 $T=39640 17490 0 0 $X=39560 $Y=17240
X127 28 M2_M1_CDNS_9 $T=43850 8260 0 0 $X=43770 $Y=8010
X128 29 M2_M1_CDNS_9 $T=43880 660 0 0 $X=43800 $Y=410
X129 30 M5_M4_CDNS_10 $T=28820 19250 0 0 $X=28740 $Y=19120
X130 33 M5_M4_CDNS_10 $T=35550 19590 0 0 $X=35470 $Y=19460
X131 1 M3_M2_CDNS_11 $T=1390 19500 0 0 $X=1310 $Y=19250
X132 21 M3_M2_CDNS_11 $T=3370 8280 0 0 $X=3290 $Y=8030
X133 43 M3_M2_CDNS_11 $T=5400 9800 0 0 $X=5320 $Y=9550
X134 7 M3_M2_CDNS_11 $T=7950 19550 0 0 $X=7870 $Y=19300
X135 25 M3_M2_CDNS_11 $T=12950 9830 0 0 $X=12870 $Y=9580
X136 44 M3_M2_CDNS_11 $T=14070 2580 0 90 $X=13820 $Y=2500
X137 39 M3_M2_CDNS_11 $T=15700 9710 0 0 $X=15620 $Y=9460
X138 11 M3_M2_CDNS_11 $T=25590 19380 0 0 $X=25510 $Y=19130
X139 35 M3_M2_CDNS_11 $T=25970 20660 0 0 $X=25890 $Y=20410
X140 46 M3_M2_CDNS_11 $T=28540 8430 0 0 $X=28460 $Y=8180
X141 46 M3_M2_CDNS_11 $T=28700 9810 0 0 $X=28620 $Y=9560
X142 32 M3_M2_CDNS_11 $T=38260 18710 0 0 $X=38180 $Y=18460
X143 42 M3_M2_CDNS_11 $T=42090 2930 0 90 $X=41840 $Y=2850
X144 1 M4_M3_CDNS_12 $T=1390 19500 0 0 $X=1310 $Y=19250
X145 21 M4_M3_CDNS_12 $T=3370 8280 0 0 $X=3290 $Y=8030
X146 7 M4_M3_CDNS_12 $T=4510 16920 0 0 $X=4430 $Y=16670
X147 43 M4_M3_CDNS_12 $T=5400 9800 0 0 $X=5320 $Y=9550
X148 7 M4_M3_CDNS_12 $T=7950 19550 0 0 $X=7870 $Y=19300
X149 36 M4_M3_CDNS_12 $T=8750 8160 0 0 $X=8670 $Y=7910
X150 37 M4_M3_CDNS_12 $T=10750 19470 0 0 $X=10670 $Y=19220
X151 38 M4_M3_CDNS_12 $T=11680 11800 0 0 $X=11600 $Y=11550
X152 25 M4_M3_CDNS_12 $T=12950 9830 0 0 $X=12870 $Y=9580
X153 11 M4_M3_CDNS_12 $T=13290 16990 0 0 $X=13210 $Y=16740
X154 44 M4_M3_CDNS_12 $T=14070 2580 0 90 $X=13820 $Y=2500
X155 39 M4_M3_CDNS_12 $T=15700 9710 0 0 $X=15620 $Y=9460
X156 38 M4_M3_CDNS_12 $T=22150 6400 0 0 $X=22070 $Y=6150
X157 39 M4_M3_CDNS_12 $T=24490 750 0 0 $X=24410 $Y=500
X158 11 M4_M3_CDNS_12 $T=25590 19380 0 0 $X=25510 $Y=19130
X159 35 M4_M3_CDNS_12 $T=25970 20660 0 0 $X=25890 $Y=20410
X160 40 M4_M3_CDNS_12 $T=26370 19410 0 0 $X=26290 $Y=19160
X161 33 M4_M3_CDNS_12 $T=26600 23000 0 0 $X=26520 $Y=22750
X162 46 M4_M3_CDNS_12 $T=28540 8430 0 0 $X=28460 $Y=8180
X163 46 M4_M3_CDNS_12 $T=28700 9810 0 0 $X=28620 $Y=9560
X164 41 M4_M3_CDNS_12 $T=29280 19170 0 0 $X=29200 $Y=18920
X165 42 M4_M3_CDNS_12 $T=35970 2380 0 0 $X=35890 $Y=2130
X166 32 M4_M3_CDNS_12 $T=38260 18710 0 0 $X=38180 $Y=18460
X167 41 M4_M3_CDNS_12 $T=39640 17490 0 0 $X=39560 $Y=17240
X168 42 M4_M3_CDNS_12 $T=42090 2930 0 90 $X=41840 $Y=2850
X169 28 M4_M3_CDNS_12 $T=43850 8260 0 0 $X=43770 $Y=8010
X170 29 M4_M3_CDNS_12 $T=43880 660 0 0 $X=43800 $Y=410
X171 32 M4_M3_CDNS_12 $T=46340 18970 0 0 $X=46260 $Y=18720
X172 1 M4_M3_CDNS_13 $T=1390 21140 0 0 $X=1310 $Y=21010
X173 21 M4_M3_CDNS_13 $T=3650 6110 0 0 $X=3570 $Y=5980
X174 43 M4_M3_CDNS_13 $T=6680 2460 0 0 $X=6600 $Y=2330
X175 35 M4_M3_CDNS_13 $T=13170 22790 0 0 $X=13090 $Y=22660
X176 25 M4_M3_CDNS_13 $T=13680 4950 0 0 $X=13600 $Y=4820
X177 11 M4_M3_CDNS_13 $T=14530 13310 0 0 $X=14450 $Y=13180
X178 11 M4_M3_CDNS_13 $T=14530 15600 0 0 $X=14450 $Y=15470
X179 44 M4_M3_CDNS_13 $T=21870 1570 0 0 $X=21790 $Y=1440
X180 36 M4_M3_CDNS_13 $T=23120 3950 0 0 $X=23040 $Y=3820
X181 40 M4_M3_CDNS_13 $T=28320 12210 0 0 $X=28240 $Y=12080
X182 29 M4_M3_CDNS_13 $T=28540 230 0 90 $X=28410 $Y=150
X183 28 M4_M3_CDNS_13 $T=28550 7610 0 90 $X=28420 $Y=7530
X184 37 M4_M3_CDNS_13 $T=33860 19960 0 90 $X=33730 $Y=19880
X185 1 M1_PO_CDNS_14 $T=1350 15570 0 0 $X=1250 $Y=15320
X186 1 M1_PO_CDNS_14 $T=1360 13320 0 0 $X=1260 $Y=13070
X187 7 M1_PO_CDNS_14 $T=4510 16920 0 0 $X=4410 $Y=16670
X188 7 M1_PO_CDNS_14 $T=5740 15570 0 0 $X=5640 $Y=15320
X189 7 M1_PO_CDNS_14 $T=5750 13320 0 0 $X=5650 $Y=13070
X190 19 M1_PO_CDNS_14 $T=6590 5910 0 0 $X=6490 $Y=5660
X191 23 M1_PO_CDNS_14 $T=7520 22860 0 0 $X=7420 $Y=22610
X192 23 M1_PO_CDNS_14 $T=7960 21030 0 0 $X=7860 $Y=20780
X193 8 M1_PO_CDNS_14 $T=8980 17010 0 0 $X=8880 $Y=16760
X194 8 M1_PO_CDNS_14 $T=10140 15570 0 0 $X=10040 $Y=15320
X195 8 M1_PO_CDNS_14 $T=10150 13320 0 0 $X=10050 $Y=13070
X196 8 M1_PO_CDNS_14 $T=10370 18740 0 0 $X=10270 $Y=18490
X197 37 M1_PO_CDNS_14 $T=10750 19470 0 0 $X=10650 $Y=19220
X198 20 M1_PO_CDNS_14 $T=12260 20780 0 0 $X=12160 $Y=20530
X199 11 M1_PO_CDNS_14 $T=13290 16990 0 0 $X=13190 $Y=16740
X200 11 M1_PO_CDNS_14 $T=14530 13310 0 0 $X=14430 $Y=13060
X201 11 M1_PO_CDNS_14 $T=14530 15600 0 0 $X=14430 $Y=15350
X202 27 M1_PO_CDNS_14 $T=14690 20780 0 0 $X=14590 $Y=20530
X203 28 M1_PO_CDNS_14 $T=15670 8330 0 0 $X=15570 $Y=8080
X204 29 M1_PO_CDNS_14 $T=16600 750 0 0 $X=16500 $Y=500
X205 38 M1_PO_CDNS_14 $T=22150 6400 0 0 $X=22050 $Y=6150
X206 39 M1_PO_CDNS_14 $T=24490 750 0 0 $X=24390 $Y=500
X207 41 M1_PO_CDNS_14 $T=29280 19170 0 0 $X=29180 $Y=18920
X208 30 M1_PO_CDNS_14 $T=34220 19150 0 0 $X=34120 $Y=18900
X209 31 M1_PO_CDNS_14 $T=35760 21100 0 0 $X=35660 $Y=20850
X210 42 M1_PO_CDNS_14 $T=35970 2380 0 0 $X=35870 $Y=2130
X211 1 M1_PO_CDNS_15 $T=1390 17230 0 0 $X=1290 $Y=16980
X212 1 M1_PO_CDNS_15 $T=1390 24660 0 0 $X=1290 $Y=24410
X213 3 M1_PO_CDNS_15 $T=2770 22320 0 90 $X=2520 $Y=22220
X214 5 M1_PO_CDNS_15 $T=2650 13610 0 0 $X=2550 $Y=13360
X215 4 M1_PO_CDNS_15 $T=2750 17050 0 0 $X=2650 $Y=16800
X216 1 M1_PO_CDNS_15 $T=4410 23850 0 0 $X=4310 $Y=23600
X217 4 M1_PO_CDNS_15 $T=5790 16970 0 0 $X=5690 $Y=16720
X218 9 M1_PO_CDNS_15 $T=7290 23970 0 90 $X=7040 $Y=23870
X219 5 M1_PO_CDNS_15 $T=7180 13450 0 0 $X=7080 $Y=13200
X220 3 M1_PO_CDNS_15 $T=8720 22330 0 90 $X=8470 $Y=22230
X221 3 M1_PO_CDNS_15 $T=9910 24890 0 90 $X=9660 $Y=24790
X222 4 M1_PO_CDNS_15 $T=10210 17010 0 0 $X=10110 $Y=16760
X223 7 M1_PO_CDNS_15 $T=11550 22710 0 0 $X=11450 $Y=22460
X224 5 M1_PO_CDNS_15 $T=11730 13390 0 0 $X=11630 $Y=13140
X225 9 M1_PO_CDNS_15 $T=13230 23970 0 90 $X=12980 $Y=23870
X226 4 M1_PO_CDNS_15 $T=14630 17040 0 0 $X=14530 $Y=16790
X227 7 M1_PO_CDNS_15 $T=15790 22330 0 90 $X=15540 $Y=22230
X228 5 M1_PO_CDNS_15 $T=15980 13520 0 0 $X=15880 $Y=13270
X229 3 M1_PO_CDNS_15 $T=17780 24480 0 0 $X=17680 $Y=24230
X230 8 M1_PO_CDNS_15 $T=20560 22320 0 90 $X=20310 $Y=22220
X231 9 M1_PO_CDNS_15 $T=22240 23950 0 0 $X=22140 $Y=23700
X232 8 M1_PO_CDNS_15 $T=24880 22320 0 90 $X=24630 $Y=22220
X233 3 M1_PO_CDNS_15 $T=26710 24400 0 0 $X=26610 $Y=24150
X234 46 M1_PO_CDNS_15 $T=28540 6330 0 0 $X=28440 $Y=6080
X235 11 M1_PO_CDNS_15 $T=29350 22530 0 0 $X=29250 $Y=22280
X236 45 M1_PO_CDNS_15 $T=29800 13490 0 0 $X=29700 $Y=13240
X237 9 M1_PO_CDNS_15 $T=31140 23850 0 0 $X=31040 $Y=23600
X238 47 M1_PO_CDNS_15 $T=31170 13680 0 0 $X=31070 $Y=13430
X239 32 M1_PO_CDNS_15 $T=31860 16950 0 0 $X=31760 $Y=16700
X240 11 M1_PO_CDNS_15 $T=33650 22300 0 90 $X=33400 $Y=22200
X241 49 M1_PO_CDNS_15 $T=35890 9730 0 0 $X=35790 $Y=9480
X242 1 M2_M1_CDNS_17 $T=1390 17230 0 0 $X=1310 $Y=16980
X243 1 M2_M1_CDNS_17 $T=1390 24660 0 0 $X=1310 $Y=24410
X244 3 M2_M1_CDNS_17 $T=2770 22320 0 90 $X=2520 $Y=22240
X245 5 M2_M1_CDNS_17 $T=2650 13610 0 0 $X=2570 $Y=13360
X246 4 M2_M1_CDNS_17 $T=2750 17050 0 0 $X=2670 $Y=16800
X247 1 M2_M1_CDNS_17 $T=4410 23850 0 0 $X=4330 $Y=23600
X248 4 M2_M1_CDNS_17 $T=5790 16970 0 0 $X=5710 $Y=16720
X249 9 M2_M1_CDNS_17 $T=7290 23970 0 90 $X=7040 $Y=23890
X250 5 M2_M1_CDNS_17 $T=7180 13450 0 0 $X=7100 $Y=13200
X251 3 M2_M1_CDNS_17 $T=8720 22330 0 90 $X=8470 $Y=22250
X252 3 M2_M1_CDNS_17 $T=9910 24890 0 90 $X=9660 $Y=24810
X253 4 M2_M1_CDNS_17 $T=10210 17010 0 0 $X=10130 $Y=16760
X254 7 M2_M1_CDNS_17 $T=11550 22710 0 0 $X=11470 $Y=22460
X255 5 M2_M1_CDNS_17 $T=11730 13390 0 0 $X=11650 $Y=13140
X256 9 M2_M1_CDNS_17 $T=13230 23970 0 90 $X=12980 $Y=23890
X257 4 M2_M1_CDNS_17 $T=14630 17040 0 0 $X=14550 $Y=16790
X258 7 M2_M1_CDNS_17 $T=15790 22330 0 90 $X=15540 $Y=22250
X259 5 M2_M1_CDNS_17 $T=15980 13520 0 0 $X=15900 $Y=13270
X260 3 M2_M1_CDNS_17 $T=17780 24480 0 0 $X=17700 $Y=24230
X261 8 M2_M1_CDNS_17 $T=20560 22320 0 90 $X=20310 $Y=22240
X262 9 M2_M1_CDNS_17 $T=22240 23950 0 0 $X=22160 $Y=23700
X263 8 M2_M1_CDNS_17 $T=24880 22320 0 90 $X=24630 $Y=22240
X264 3 M2_M1_CDNS_17 $T=26710 24400 0 0 $X=26630 $Y=24150
X265 46 M2_M1_CDNS_17 $T=28540 6330 0 0 $X=28460 $Y=6080
X266 11 M2_M1_CDNS_17 $T=29350 22530 0 0 $X=29270 $Y=22280
X267 45 M2_M1_CDNS_17 $T=29800 13490 0 0 $X=29720 $Y=13240
X268 9 M2_M1_CDNS_17 $T=31140 23850 0 0 $X=31060 $Y=23600
X269 47 M2_M1_CDNS_17 $T=31170 13680 0 0 $X=31090 $Y=13430
X270 32 M2_M1_CDNS_17 $T=31860 16950 0 0 $X=31780 $Y=16700
X271 11 M2_M1_CDNS_17 $T=33650 22300 0 90 $X=33400 $Y=22220
X272 49 M2_M1_CDNS_17 $T=35890 9730 0 0 $X=35810 $Y=9480
X273 1 6 2 5 43 77 AND $T=40 14460 1 0 $X=50 $Y=10660
X274 1 6 2 4 21 76 AND $T=40 14420 0 0 $X=50 $Y=14420
X275 1 6 2 3 20 75 AND $T=40 21740 0 0 $X=50 $Y=21740
X276 7 6 2 5 39 80 AND $T=4440 14460 1 0 $X=4450 $Y=10660
X277 7 6 2 4 24 79 AND $T=4440 14420 0 0 $X=4450 $Y=14420
X278 1 6 2 9 23 78 AND $T=4440 21740 0 0 $X=4450 $Y=21740
X279 8 6 2 5 38 83 AND $T=8840 14460 1 0 $X=8850 $Y=10660
X280 8 6 2 4 26 82 AND $T=8840 14420 0 0 $X=8850 $Y=14420
X281 3 6 2 7 35 81 AND $T=8840 21740 0 0 $X=8850 $Y=21740
X282 11 6 2 5 50 93 AND $T=13240 14460 1 0 $X=13250 $Y=10660
X283 11 6 2 4 45 92 AND $T=13240 14420 0 0 $X=13250 $Y=14420
X284 9 6 2 7 27 91 AND $T=13240 21740 0 0 $X=13250 $Y=21740
X285 3 6 2 8 30 104 AND $T=17880 21740 0 0 $X=17890 $Y=21740
X286 9 6 2 8 33 126 AND $T=22280 21740 0 0 $X=22290 $Y=21740
X287 3 6 2 11 14 127 AND $T=26680 21740 0 0 $X=26690 $Y=21740
X288 9 6 2 11 31 131 AND $T=31080 21740 0 0 $X=31090 $Y=21740
X289 23 2 6 37 22 25 73 74 225 half_adder $T=50 21780 1 0 $X=50 $Y=17980
X290 50 2 6 48 13 46 102 103 228 half_adder $T=17640 14460 1 0 $X=17640 $Y=10660
X291 45 2 6 47 17 49 129 130 237 half_adder $T=29830 14460 1 0 $X=29830 $Y=10660
X292 30 2 6 31 18 32 133 134 238 half_adder $T=34210 21780 1 0 $X=34210 $Y=17980
X293 22 6 24 2 28 36 19 67 70 71
+ 65 66 68 69 223 224 full_adder1_small $T=22270 7090 1 180 $X=20 $Y=7100
X294 43 6 34 2 29 10 12 60 63 64
+ 58 59 61 62 221 222 full_adder1_small $T=30 -230 0 0 $X=50 $Y=-220
X295 21 6 25 2 19 44 34 53 56 57
+ 51 52 54 55 219 220 full_adder1_small $T=30 7150 1 0 $X=50 $Y=3340
X296 20 6 27 2 41 40 37 86 89 90
+ 84 85 87 88 226 227 full_adder1_small $T=12230 21790 1 0 $X=12250 $Y=17980
X297 33 6 35 2 32 47 41 96 99 100
+ 94 95 97 98 229 230 full_adder1_small $T=17850 14410 0 0 $X=17870 $Y=14420
X298 39 6 44 2 42 15 29 121 124 125
+ 119 120 122 123 235 236 full_adder1_small $T=21990 -230 0 0 $X=22010 $Y=-220
X299 38 6 36 2 46 16 42 114 117 118
+ 112 113 115 116 233 234 full_adder1_small $T=21990 7150 1 0 $X=22010 $Y=3340
X300 26 6 40 2 49 48 28 107 110 111
+ 105 106 108 109 231 232 full_adder1_small $T=21990 7090 0 0 $X=22010 $Y=7100
M0 77 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=11610 $dt=1
M1 76 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=16790 $dt=1
M2 75 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5317 scb=0.0167655 scc=0.000436143 $X=740 $Y=24110 $dt=1
M3 73 23 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=16.2188 scb=0.0173423 scc=0.000698846 $X=750 $Y=18640 $dt=1
M4 58 43 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=2120 $dt=1
M5 51 21 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=820 $Y=4320 $dt=1
M6 19 71 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=1070 $Y=9450 $dt=1
M7 6 70 19 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=1480 $Y=9450 $dt=1
M8 59 34 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=2120 $dt=1
M9 52 25 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1780 $Y=4320 $dt=1
M10 77 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=11600 $dt=1
M11 76 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=16800 $dt=1
M12 75 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.96224 scb=0.0072004 scc=0.000178239 $X=1980 $Y=24120 $dt=1
M13 221 34 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=1880 $dt=1
M14 219 25 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3110 $Y=4080 $dt=1
M15 43 77 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=11580 $dt=1
M16 21 76 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=16820 $dt=1
M17 20 75 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=3660 $Y=24140 $dt=1
M18 71 24 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=3910 $Y=9450 $dt=1
M19 60 58 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=1940 $dt=1
M20 53 51 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4080 $Y=4020 $dt=1
M21 6 22 71 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=4320 $Y=9450 $dt=1
M22 60 59 221 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=1940 $dt=1
M23 53 52 219 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5040 $Y=4020 $dt=1
M24 80 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=11610 $dt=1
M25 79 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=16790 $dt=1
M26 78 1 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5140 $Y=24110 $dt=1
M27 221 43 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=1940 $dt=1
M28 219 21 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6000 $Y=4020 $dt=1
M29 22 37 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=6190 $Y=18700 $dt=1
M30 80 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=11600 $dt=1
M31 79 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=16800 $dt=1
M32 78 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6380 $Y=24120 $dt=1
M33 70 67 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=6890 $Y=9230 $dt=1
M34 6 28 70 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=7300 $Y=9230 $dt=1
M35 22 23 225 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=7300 $Y=18660 $dt=1
M36 61 29 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=2120 $dt=1
M37 54 19 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7660 $Y=4320 $dt=1
M38 39 80 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=11580 $dt=1
M39 24 79 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=16820 $dt=1
M40 23 78 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=8060 $Y=24140 $dt=1
M41 74 23 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=8540 $Y=18930 $dt=1
M42 62 60 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=2120 $dt=1
M43 55 53 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8620 $Y=4320 $dt=1
M44 6 28 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=9370 $Y=9260 $dt=1
M45 83 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=11610 $dt=1
M46 82 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=16790 $dt=1
M47 81 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=9540 $Y=24110 $dt=1
M48 74 37 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=9780 $Y=18920 $dt=1
M49 222 60 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=1880 $dt=1
M50 220 53 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9950 $Y=4080 $dt=1
M51 224 69 36 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10330 $Y=9260 $dt=1
M52 83 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=11600 $dt=1
M53 82 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=16800 $dt=1
M54 81 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=10780 $Y=24120 $dt=1
M55 10 61 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=1940 $dt=1
M56 44 54 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10920 $Y=4020 $dt=1
M57 224 68 36 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11290 $Y=9260 $dt=1
M58 25 74 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=11460 $Y=18900 $dt=1
M59 10 62 222 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=1940 $dt=1
M60 44 55 220 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11880 $Y=4020 $dt=1
M61 6 67 224 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=12260 $Y=9200 $dt=1
M62 38 83 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=11580 $dt=1
M63 26 82 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=16820 $dt=1
M64 35 81 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=12460 $Y=24140 $dt=1
M65 222 29 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=1940 $dt=1
M66 220 19 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12840 $Y=4020 $dt=1
M67 84 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13020 $Y=18960 $dt=1
M68 6 67 69 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13590 $Y=9440 $dt=1
M69 93 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=11610 $dt=1
M70 92 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=16790 $dt=1
M71 91 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=13940 $Y=24110 $dt=1
M72 85 27 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=13980 $Y=18960 $dt=1
M73 6 28 68 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=14550 $Y=9440 $dt=1
M74 63 29 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=1910 $dt=1
M75 56 19 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14910 $Y=4050 $dt=1
M76 93 5 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=11600 $dt=1
M77 92 4 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=16800 $dt=1
M78 91 7 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=15180 $Y=24120 $dt=1
M79 226 27 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=15310 $Y=18720 $dt=1
M80 6 60 63 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=1910 $dt=1
M81 6 53 56 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15320 $Y=4050 $dt=1
M82 6 22 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16210 $Y=9260 $dt=1
M83 86 84 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=16280 $Y=18660 $dt=1
M84 50 93 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=11580 $dt=1
M85 45 92 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=16820 $dt=1
M86 27 91 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=16860 $Y=24140 $dt=1
M87 223 66 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17170 $Y=9260 $dt=1
M88 86 85 226 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=17240 $Y=18660 $dt=1
M89 64 43 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=2130 $dt=1
M90 57 21 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17890 $Y=4310 $dt=1
M91 223 65 67 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18130 $Y=9260 $dt=1
M92 226 20 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=18200 $Y=18660 $dt=1
M93 6 34 64 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=2130 $dt=1
M94 6 25 57 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18300 $Y=4310 $dt=1
M95 102 50 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=18340 $Y=11320 $dt=1
M96 104 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=18580 $Y=24110 $dt=1
M97 94 33 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=18640 $Y=16760 $dt=1
M98 6 24 223 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=19100 $Y=9200 $dt=1
M99 95 35 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19600 $Y=16760 $dt=1
M100 104 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=19820 $Y=24120 $dt=1
M101 87 41 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=19860 $Y=18960 $dt=1
M102 6 24 66 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20430 $Y=9440 $dt=1
M103 12 63 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=2130 $dt=1
M104 34 56 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=20730 $Y=4310 $dt=1
M105 88 86 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=20820 $Y=18960 $dt=1
M106 229 35 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=20930 $Y=16520 $dt=1
M107 6 64 12 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=2130 $dt=1
M108 6 57 34 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21140 $Y=4310 $dt=1
M109 6 22 65 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=21390 $Y=9440 $dt=1
M110 30 104 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=21500 $Y=24140 $dt=1
M111 96 94 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=21900 $Y=16580 $dt=1
M112 227 86 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=22150 $Y=18720 $dt=1
M113 119 39 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=2120 $dt=1
M114 112 38 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=4320 $dt=1
M115 105 26 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=22780 $Y=9440 $dt=1
M116 96 95 229 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=22860 $Y=16580 $dt=1
M117 126 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=22980 $Y=24110 $dt=1
M118 40 87 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23120 $Y=18660 $dt=1
M119 120 44 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=2120 $dt=1
M120 113 36 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=4320 $dt=1
M121 106 40 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23740 $Y=9440 $dt=1
M122 13 48 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=23780 $Y=11380 $dt=1
M123 229 33 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=23820 $Y=16580 $dt=1
M124 40 88 227 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24080 $Y=18660 $dt=1
M125 126 8 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=24220 $Y=24120 $dt=1
M126 13 50 228 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=24890 $Y=11340 $dt=1
M127 227 41 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=25040 $Y=18660 $dt=1
M128 235 44 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=1880 $dt=1
M129 233 36 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=4080 $dt=1
M130 231 40 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25070 $Y=9200 $dt=1
M131 97 32 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=25480 $Y=16760 $dt=1
M132 33 126 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=25900 $Y=24140 $dt=1
M133 121 119 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=1940 $dt=1
M134 114 112 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=4020 $dt=1
M135 107 105 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26040 $Y=9260 $dt=1
M136 103 50 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26130 $Y=11610 $dt=1
M137 98 96 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=26440 $Y=16760 $dt=1
M138 121 120 235 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=1940 $dt=1
M139 114 113 233 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=4020 $dt=1
M140 107 106 231 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27000 $Y=9260 $dt=1
M141 89 41 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27110 $Y=18690 $dt=1
M142 103 48 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27370 $Y=11600 $dt=1
M143 127 3 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=27380 $Y=24110 $dt=1
M144 6 86 89 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=27520 $Y=18690 $dt=1
M145 230 96 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=27770 $Y=16520 $dt=1
M146 235 39 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=1940 $dt=1
M147 233 38 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=4020 $dt=1
M148 231 26 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27960 $Y=9260 $dt=1
M149 127 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=28620 $Y=24120 $dt=1
M150 47 97 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28740 $Y=16580 $dt=1
M151 46 103 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=29050 $Y=11580 $dt=1
M152 122 42 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=2120 $dt=1
M153 115 46 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=4320 $dt=1
M154 108 49 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=29620 $Y=9440 $dt=1
M155 47 98 230 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=29700 $Y=16580 $dt=1
M156 90 20 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30090 $Y=18950 $dt=1
M157 14 127 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.58543 scb=0.00668222 scc=0.000150123 $X=30300 $Y=24140 $dt=1
M158 6 27 90 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=30500 $Y=18950 $dt=1
M159 129 45 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=30530 $Y=11320 $dt=1
M160 123 121 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=2120 $dt=1
M161 116 114 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=4320 $dt=1
M162 109 107 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30580 $Y=9440 $dt=1
M163 230 32 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=30660 $Y=16580 $dt=1
M164 131 9 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=31780 $Y=24110 $dt=1
M165 236 121 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=1880 $dt=1
M166 234 114 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=4080 $dt=1
M167 232 107 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=31910 $Y=9200 $dt=1
M168 99 32 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=32730 $Y=16550 $dt=1
M169 15 122 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=1940 $dt=1
M170 16 115 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=4020 $dt=1
M171 48 108 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=32880 $Y=9260 $dt=1
M172 37 89 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=32930 $Y=18950 $dt=1
M173 131 11 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=33020 $Y=24120 $dt=1
M174 6 96 99 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=33140 $Y=16550 $dt=1
M175 6 90 37 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=33340 $Y=18950 $dt=1
M176 15 123 236 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=1940 $dt=1
M177 16 116 234 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=4020 $dt=1
M178 48 109 232 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33840 $Y=9260 $dt=1
M179 31 131 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=34700 $Y=24140 $dt=1
M180 236 42 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=1940 $dt=1
M181 234 46 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=4020 $dt=1
M182 232 49 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34800 $Y=9260 $dt=1
M183 133 30 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=9.94249 scb=0.00836239 scc=0.000476878 $X=34910 $Y=18640 $dt=1
M184 100 33 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=35710 $Y=16770 $dt=1
M185 17 47 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=11.6393 scb=0.010126 scc=0.000764642 $X=35970 $Y=11380 $dt=1
M186 6 35 100 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=36120 $Y=16770 $dt=1
M187 124 42 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=1910 $dt=1
M188 117 46 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=4050 $dt=1
M189 110 49 6 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=36870 $Y=9230 $dt=1
M190 17 45 237 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=37080 $Y=11340 $dt=1
M191 6 121 124 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=1910 $dt=1
M192 6 114 117 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=4050 $dt=1
M193 6 107 110 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37280 $Y=9230 $dt=1
M194 130 45 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=38320 $Y=11610 $dt=1
M195 41 99 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=38550 $Y=16770 $dt=1
M196 6 100 41 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=38960 $Y=16770 $dt=1
M197 130 47 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=39560 $Y=11600 $dt=1
M198 125 39 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=2130 $dt=1
M199 118 38 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=4310 $dt=1
M200 111 26 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=39850 $Y=9450 $dt=1
M201 6 44 125 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=2130 $dt=1
M202 6 36 118 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=4310 $dt=1
M203 6 40 111 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40260 $Y=9450 $dt=1
M204 18 31 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.2705 scb=0.0126902 scc=0.000796523 $X=40350 $Y=18700 $dt=1
M205 49 130 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7599 scb=0.0102397 scc=0.000176803 $X=41240 $Y=11580 $dt=1
M206 18 30 238 6 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=41460 $Y=18660 $dt=1
M207 29 124 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=2130 $dt=1
M208 42 117 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=42690 $Y=4310 $dt=1
M209 28 110 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=42690 $Y=9450 $dt=1
M210 134 30 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42700 $Y=18930 $dt=1
M211 6 125 29 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=2130 $dt=1
M212 6 118 42 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=43100 $Y=4310 $dt=1
M213 6 111 28 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=43100 $Y=9450 $dt=1
M214 134 31 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43940 $Y=18920 $dt=1
M215 32 134 6 6 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.8846 scb=0.00870518 scc=0.000160728 $X=45620 $Y=18900 $dt=1
.ends multiplier

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_31                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_31 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_31

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nmos1v_CDNS_32                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nmos1v_CDNS_32 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=0
.ends nmos1v_CDNS_32

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_43                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_43 1 2 3 5 6 8
*.DEVICECLIMB
** N=14 EP=6 FDC=2
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.04018 scb=0.00737277 scc=0.00014625 $X=810 $Y=710 $dt=0
M1 8 6 2 2 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.22651 scb=0.00772413 scc=0.000211444 $X=4640 $Y=580 $dt=0
.ends cellTmpl_CDNS_43

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_44                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_44 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_44

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pmos1v_CDNS_45                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pmos1v_CDNS_45 1 2 3 4 5
*.DEVICECLIMB
** N=5 EP=5 FDC=0
.ends pmos1v_CDNS_45

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X                                   *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X 1 2 3 4 5 6 7 8 9 10
+ 11 12
** N=12 EP=12 FDC=12
X0 7 M3_M2_CDNS_1 $T=250 -3000 0 0 $X=170 $Y=-3250
X1 7 M3_M2_CDNS_1 $T=960 -2040 0 0 $X=880 $Y=-2290
X2 7 M3_M2_CDNS_1 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X3 7 M2_M1_CDNS_2 $T=960 -2040 0 0 $X=880 $Y=-2290
X4 7 M2_M1_CDNS_9 $T=250 -3000 0 0 $X=170 $Y=-3250
X5 7 M2_M1_CDNS_9 $T=2620 -2730 0 0 $X=2540 $Y=-2980
X6 7 M1_PO_CDNS_14 $T=250 -3000 0 0 $X=150 $Y=-3250
X7 7 M1_PO_CDNS_14 $T=2620 -2730 0 0 $X=2520 $Y=-2980
X8 1 M1_PO_CDNS_15 $T=1300 -3500 0 0 $X=1200 $Y=-3750
X9 1 M1_PO_CDNS_15 $T=2660 -4240 0 0 $X=2560 $Y=-4490
X10 1 M1_PO_CDNS_16 $T=680 -3550 0 0 $X=580 $Y=-3670
X11 2 M1_PO_CDNS_16 $T=1300 -2090 0 0 $X=1200 $Y=-2210
X12 5 M1_PO_CDNS_16 $T=4040 -3180 0 0 $X=3940 $Y=-3300
X13 8 M1_PO_CDNS_16 $T=4300 -3670 0 90 $X=4180 $Y=-3770
X14 1 M2_M1_CDNS_17 $T=1300 -3500 0 0 $X=1220 $Y=-3750
X15 1 M2_M1_CDNS_17 $T=2660 -4240 0 0 $X=2580 $Y=-4490
X16 4 7 9 4 nmos1v_CDNS_31 $T=1990 -4420 0 0 $X=1790 $Y=-4620
X17 8 5 10 4 nmos1v_CDNS_31 $T=3370 -4430 0 0 $X=3170 $Y=-4630
X18 8 2 9 4 nmos1v_CDNS_32 $T=1780 -4420 0 0 $X=1360 $Y=-4620
X19 4 1 10 4 nmos1v_CDNS_32 $T=3160 -4430 0 0 $X=2740 $Y=-4630
X20 3 4 1 7 8 6 cellTmpl_CDNS_43 $T=-60 -5080 0 0 $X=-180 $Y=-5220
X21 3 1 11 4 3 pmos1v_CDNS_44 $T=1990 -3120 0 0 $X=1790 $Y=-3320
X22 8 5 12 4 3 pmos1v_CDNS_44 $T=3370 -3190 0 0 $X=3170 $Y=-3390
X23 8 2 11 4 3 pmos1v_CDNS_45 $T=1780 -3120 0 0 $X=1360 $Y=-3320
X24 3 7 12 4 3 pmos1v_CDNS_45 $T=3160 -3190 0 0 $X=2740 $Y=-3390
M0 9 2 8 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1780 $Y=-4420 $dt=0
M1 4 7 9 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1990 $Y=-4420 $dt=0
M2 10 1 4 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3160 $Y=-4430 $dt=0
M3 8 5 10 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3370 $Y=-4430 $dt=0
M4 7 1 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=750 $Y=-2850 $dt=1
M5 11 2 8 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1780 $Y=-3120 $dt=1
M6 3 1 11 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=1990 $Y=-3120 $dt=1
M7 12 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3160 $Y=-3190 $dt=1
M8 8 5 12 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=3370 $Y=-3190 $dt=1
M9 6 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=20.2373 scb=0.0194294 scc=0.00149528 $X=4580 $Y=-3180 $dt=1
.ends MUX_2to1___2X

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: FA_4bit                                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt FA_4bit 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19
** N=83 EP=19 FDC=144
X0 17 M3_M2_CDNS_1 $T=18840 8310 0 0 $X=18760 $Y=8060
X1 17 M3_M2_CDNS_4 $T=21980 9220 0 0 $X=21900 $Y=9090
X2 18 M3_M2_CDNS_7 $T=14030 6120 0 0 $X=13950 $Y=5870
X3 19 M3_M2_CDNS_7 $T=16960 11880 0 0 $X=16880 $Y=11630
X4 19 M3_M2_CDNS_7 $T=22610 11350 0 0 $X=22530 $Y=11100
X5 5 M2_M1_CDNS_8 $T=-80 3540 0 0 $X=-160 $Y=3410
X6 5 M2_M1_CDNS_8 $T=-80 10890 0 0 $X=-160 $Y=10760
X7 18 M2_M1_CDNS_8 $T=21770 2020 0 0 $X=21690 $Y=1890
X8 17 M2_M1_CDNS_8 $T=21770 5100 0 0 $X=21690 $Y=4970
X9 18 M2_M1_CDNS_9 $T=14030 6120 0 0 $X=13950 $Y=5870
X10 19 M2_M1_CDNS_9 $T=16960 11880 0 0 $X=16880 $Y=11630
X11 17 M2_M1_CDNS_9 $T=18840 8310 0 0 $X=18760 $Y=8060
X12 19 M2_M1_CDNS_9 $T=22610 11350 0 0 $X=22530 $Y=11100
X13 18 M3_M2_CDNS_11 $T=19730 4760 0 0 $X=19650 $Y=4510
X14 18 M4_M3_CDNS_12 $T=14030 6120 0 0 $X=13950 $Y=5870
X15 19 M4_M3_CDNS_12 $T=16960 11880 0 0 $X=16880 $Y=11630
X16 18 M4_M3_CDNS_12 $T=19730 4760 0 0 $X=19650 $Y=4510
X17 19 M4_M3_CDNS_12 $T=22610 11350 0 0 $X=22530 $Y=11100
X18 18 M1_PO_CDNS_14 $T=14030 6120 0 0 $X=13930 $Y=5870
X19 19 M1_PO_CDNS_14 $T=16960 11880 0 0 $X=16860 $Y=11630
X20 17 M1_PO_CDNS_14 $T=18840 8310 0 0 $X=18740 $Y=8060
X21 6 5 1 7 11 12 18 43 46 47
+ 41 42 44 45 82 83 full_adder1_small $T=-90 -130 0 0 $X=-70 $Y=-120
X22 8 5 2 7 18 13 17 36 39 40
+ 34 35 37 38 80 81 full_adder1_small $T=-90 7250 1 0 $X=-70 $Y=3440
X23 9 5 3 7 17 14 19 29 32 33
+ 27 28 30 31 78 79 full_adder1_small $T=-90 7190 0 0 $X=-70 $Y=7200
X24 10 5 4 7 19 15 16 22 25 26
+ 20 21 23 24 76 77 full_adder1_small $T=-90 14570 1 0 $X=-70 $Y=10760
M0 41 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=2220 $dt=1
M1 34 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=4420 $dt=1
M2 27 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=9540 $dt=1
M3 20 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.672 scb=0.0152131 scc=0.000371293 $X=700 $Y=11740 $dt=1
M4 42 1 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=2220 $dt=1
M5 35 2 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=4420 $dt=1
M6 28 3 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=9540 $dt=1
M7 21 4 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=1660 $Y=11740 $dt=1
M8 82 1 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=1980 $dt=1
M9 80 2 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=4180 $dt=1
M10 78 3 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=9300 $dt=1
M11 76 4 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=2990 $Y=11500 $dt=1
M12 43 41 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=2040 $dt=1
M13 36 34 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=4120 $dt=1
M14 29 27 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=9360 $dt=1
M15 22 20 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=3960 $Y=11440 $dt=1
M16 43 42 82 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=2040 $dt=1
M17 36 35 80 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=4120 $dt=1
M18 29 28 78 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=9360 $dt=1
M19 22 21 76 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4920 $Y=11440 $dt=1
M20 82 6 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=2040 $dt=1
M21 80 8 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=4120 $dt=1
M22 78 9 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=9360 $dt=1
M23 76 10 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5880 $Y=11440 $dt=1
M24 44 11 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=2220 $dt=1
M25 37 18 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=4420 $dt=1
M26 30 17 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=9540 $dt=1
M27 23 19 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=7540 $Y=11740 $dt=1
M28 45 43 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=2220 $dt=1
M29 38 36 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=4420 $dt=1
M30 31 29 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=9540 $dt=1
M31 24 22 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8500 $Y=11740 $dt=1
M32 83 43 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=1980 $dt=1
M33 81 36 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=4180 $dt=1
M34 79 29 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=9300 $dt=1
M35 77 22 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=9830 $Y=11500 $dt=1
M36 12 44 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=2040 $dt=1
M37 13 37 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=4120 $dt=1
M38 14 30 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=9360 $dt=1
M39 15 23 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=10800 $Y=11440 $dt=1
M40 12 45 83 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=2040 $dt=1
M41 13 38 81 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=4120 $dt=1
M42 14 31 79 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=9360 $dt=1
M43 15 24 77 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11760 $Y=11440 $dt=1
M44 83 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=2040 $dt=1
M45 81 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=4120 $dt=1
M46 79 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=9360 $dt=1
M47 77 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12720 $Y=11440 $dt=1
M48 46 11 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=2010 $dt=1
M49 39 18 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=4150 $dt=1
M50 32 17 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=9330 $dt=1
M51 25 19 5 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=14790 $Y=11470 $dt=1
M52 5 43 46 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=2010 $dt=1
M53 5 36 39 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=4150 $dt=1
M54 5 29 32 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=9330 $dt=1
M55 5 22 25 5 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15200 $Y=11470 $dt=1
M56 47 6 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=2230 $dt=1
M57 40 8 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=4410 $dt=1
M58 33 9 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=9550 $dt=1
M59 26 10 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=17770 $Y=11730 $dt=1
M60 5 1 47 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=2230 $dt=1
M61 5 2 40 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=4410 $dt=1
M62 5 3 33 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=9550 $dt=1
M63 5 4 26 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18180 $Y=11730 $dt=1
M64 18 46 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=2230 $dt=1
M65 17 39 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=4410 $dt=1
M66 19 32 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=9550 $dt=1
M67 16 25 5 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=10.287 scb=0.00843354 scc=0.000230522 $X=20610 $Y=11730 $dt=1
M68 5 47 18 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=2230 $dt=1
M69 5 40 17 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=4410 $dt=1
M70 5 33 19 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=9550 $dt=1
M71 5 26 16 5 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.9797 scb=0.0105745 scc=0.000243193 $X=21020 $Y=11730 $dt=1
.ends FA_4bit

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small 1 2 3 4
** N=4 EP=4 FDC=2
X0 1 M1_PO_CDNS_16 $T=950 1780 0 90 $X=830 $Y=1680
X1 2 3 cellTmpl_CDNS_18 $T=120 140 0 0 $X=0 $Y=0
M0 4 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.7353 scb=0.0117274 scc=0.000445561 $X=1070 $Y=980 $dt=0
M1 4 1 2 2 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8675 scb=0.0146094 scc=0.000688105 $X=1070 $Y=2220 $dt=1
.ends INV_1X_small

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: 10badder                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt 10badder 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 64
+ 65 66 67 68 69 70 149 150 151 152
+ 153 154 155 256 257 266 267
*.DEVICECLIMB
** N=267 EP=77 FDC=483
X0 2 M3_M2_CDNS_1 $T=52330 32180 0 90 $X=52080 $Y=32100
X1 35 M3_M2_CDNS_1 $T=52330 46820 0 90 $X=52080 $Y=46740
X2 36 M3_M2_CDNS_1 $T=53480 29020 0 0 $X=53400 $Y=28770
X3 37 M3_M2_CDNS_1 $T=53480 43660 0 0 $X=53400 $Y=43410
X4 38 M3_M2_CDNS_1 $T=54270 29810 0 90 $X=54020 $Y=29730
X5 39 M3_M2_CDNS_1 $T=54270 44450 0 90 $X=54020 $Y=44370
X6 36 M3_M2_CDNS_1 $T=55540 26280 0 0 $X=55460 $Y=26030
X7 37 M3_M2_CDNS_1 $T=55540 40920 0 0 $X=55460 $Y=40670
X8 40 M3_M2_CDNS_1 $T=55730 21200 0 90 $X=55480 $Y=21120
X9 41 M3_M2_CDNS_1 $T=55730 35840 0 90 $X=55480 $Y=35760
X10 42 M3_M2_CDNS_1 $T=56210 23810 0 90 $X=55960 $Y=23730
X11 43 M3_M2_CDNS_1 $T=56210 38450 0 90 $X=55960 $Y=38370
X12 44 M3_M2_CDNS_1 $T=56050 31070 0 0 $X=55970 $Y=30820
X13 45 M3_M2_CDNS_1 $T=56050 45710 0 0 $X=55970 $Y=45460
X14 46 M3_M2_CDNS_1 $T=56240 34220 0 0 $X=56160 $Y=33970
X15 47 M3_M2_CDNS_1 $T=56240 48860 0 0 $X=56160 $Y=48610
X16 13 M3_M2_CDNS_1 $T=57660 26200 0 90 $X=57410 $Y=26120
X17 11 M3_M2_CDNS_1 $T=57660 33520 0 90 $X=57410 $Y=33440
X18 10 M3_M2_CDNS_1 $T=57660 40840 0 90 $X=57410 $Y=40760
X19 8 M3_M2_CDNS_1 $T=57660 48160 0 90 $X=57410 $Y=48080
X20 7 M3_M2_CDNS_1 $T=57670 22770 0 90 $X=57420 $Y=22690
X21 12 M3_M2_CDNS_1 $T=57670 30070 0 90 $X=57420 $Y=29990
X22 6 M3_M2_CDNS_1 $T=57670 37410 0 90 $X=57420 $Y=37330
X23 9 M3_M2_CDNS_1 $T=57670 44710 0 90 $X=57420 $Y=44630
X24 44 M3_M2_CDNS_1 $T=62950 31240 0 90 $X=62700 $Y=31160
X25 45 M3_M2_CDNS_1 $T=62950 45880 0 90 $X=62700 $Y=45800
X26 42 M3_M2_CDNS_1 $T=63400 23460 0 0 $X=63320 $Y=23210
X27 43 M3_M2_CDNS_1 $T=63400 38100 0 0 $X=63320 $Y=37850
X28 40 M3_M2_CDNS_1 $T=63720 21760 0 0 $X=63640 $Y=21510
X29 41 M3_M2_CDNS_1 $T=63720 36400 0 0 $X=63640 $Y=36150
X30 38 M3_M2_CDNS_1 $T=63820 29420 0 0 $X=63740 $Y=29170
X31 39 M3_M2_CDNS_1 $T=63820 44060 0 0 $X=63740 $Y=43810
X32 36 M2_M1_CDNS_2 $T=53480 29020 0 0 $X=53400 $Y=28770
X33 37 M2_M1_CDNS_2 $T=53480 43660 0 0 $X=53400 $Y=43410
X34 46 M2_M1_CDNS_2 $T=56240 34220 0 0 $X=56160 $Y=33970
X35 47 M2_M1_CDNS_2 $T=56240 48860 0 0 $X=56160 $Y=48610
X36 44 M2_M1_CDNS_2 $T=62950 31240 0 90 $X=62700 $Y=31160
X37 45 M2_M1_CDNS_2 $T=62950 45880 0 90 $X=62700 $Y=45800
X38 42 M2_M1_CDNS_2 $T=63400 23460 0 0 $X=63320 $Y=23210
X39 43 M2_M1_CDNS_2 $T=63400 38100 0 0 $X=63320 $Y=37850
X40 40 M2_M1_CDNS_2 $T=63720 21760 0 0 $X=63640 $Y=21510
X41 41 M2_M1_CDNS_2 $T=63720 36400 0 0 $X=63640 $Y=36150
X42 38 M2_M1_CDNS_2 $T=63820 29420 0 0 $X=63740 $Y=29170
X43 39 M2_M1_CDNS_2 $T=63820 44060 0 0 $X=63740 $Y=43810
X44 46 M3_M2_CDNS_4 $T=50730 34460 0 0 $X=50650 $Y=34330
X45 47 M3_M2_CDNS_4 $T=50800 49100 0 0 $X=50720 $Y=48970
X46 2 M3_M2_CDNS_4 $T=51610 22610 0 0 $X=51530 $Y=22480
X47 35 M3_M2_CDNS_7 $T=51080 34160 0 0 $X=51000 $Y=33910
X48 48 M3_M2_CDNS_7 $T=56340 32800 0 0 $X=56260 $Y=32550
X49 49 M3_M2_CDNS_7 $T=56340 47440 0 0 $X=56260 $Y=47190
X50 50 M3_M2_CDNS_7 $T=57240 50840 0 0 $X=57160 $Y=50590
X51 51 M3_M2_CDNS_7 $T=72650 52420 0 90 $X=72400 $Y=52340
X52 35 M3_M2_CDNS_7 $T=78550 36430 0 0 $X=78470 $Y=36180
X53 51 M3_M2_CDNS_7 $T=79400 52420 0 90 $X=79150 $Y=52340
X54 48 M3_M2_CDNS_7 $T=86760 34460 0 0 $X=86680 $Y=34210
X55 49 M3_M2_CDNS_7 $T=86760 49100 0 0 $X=86680 $Y=48850
X56 3 M2_M1_CDNS_8 $T=50480 50560 0 0 $X=50400 $Y=50430
X57 3 M2_M1_CDNS_8 $T=51590 45750 0 90 $X=51460 $Y=45670
X58 46 M2_M1_CDNS_8 $T=53210 27000 0 0 $X=53130 $Y=26870
X59 47 M2_M1_CDNS_8 $T=53210 41640 0 0 $X=53130 $Y=41510
X60 52 M2_M1_CDNS_8 $T=53230 23140 0 0 $X=53150 $Y=23010
X61 53 M2_M1_CDNS_8 $T=53230 37780 0 0 $X=53150 $Y=37650
X62 3 M2_M1_CDNS_8 $T=62920 24380 0 0 $X=62840 $Y=24250
X63 3 M2_M1_CDNS_8 $T=62920 39020 0 0 $X=62840 $Y=38890
X64 3 M2_M1_CDNS_8 $T=62930 31710 0 0 $X=62850 $Y=31580
X65 3 M2_M1_CDNS_8 $T=62930 46350 0 0 $X=62850 $Y=46220
X66 35 M2_M1_CDNS_9 $T=51080 34160 0 0 $X=51000 $Y=33910
X67 2 M2_M1_CDNS_9 $T=52330 32180 0 90 $X=52080 $Y=32100
X68 35 M2_M1_CDNS_9 $T=52330 46820 0 90 $X=52080 $Y=46740
X69 38 M2_M1_CDNS_9 $T=54270 29810 0 90 $X=54020 $Y=29730
X70 39 M2_M1_CDNS_9 $T=54270 44450 0 90 $X=54020 $Y=44370
X71 36 M2_M1_CDNS_9 $T=55540 26280 0 0 $X=55460 $Y=26030
X72 37 M2_M1_CDNS_9 $T=55540 40920 0 0 $X=55460 $Y=40670
X73 40 M2_M1_CDNS_9 $T=55730 21200 0 90 $X=55480 $Y=21120
X74 41 M2_M1_CDNS_9 $T=55730 35840 0 90 $X=55480 $Y=35760
X75 42 M2_M1_CDNS_9 $T=56210 23810 0 90 $X=55960 $Y=23730
X76 43 M2_M1_CDNS_9 $T=56210 38450 0 90 $X=55960 $Y=38370
X77 44 M2_M1_CDNS_9 $T=56050 31070 0 0 $X=55970 $Y=30820
X78 45 M2_M1_CDNS_9 $T=56050 45710 0 0 $X=55970 $Y=45460
X79 48 M2_M1_CDNS_9 $T=56340 32800 0 0 $X=56260 $Y=32550
X80 49 M2_M1_CDNS_9 $T=56340 47440 0 0 $X=56260 $Y=47190
X81 50 M2_M1_CDNS_9 $T=57240 50840 0 0 $X=57160 $Y=50590
X82 13 M2_M1_CDNS_9 $T=57660 26200 0 90 $X=57410 $Y=26120
X83 11 M2_M1_CDNS_9 $T=57660 33520 0 90 $X=57410 $Y=33440
X84 10 M2_M1_CDNS_9 $T=57660 40840 0 90 $X=57410 $Y=40760
X85 8 M2_M1_CDNS_9 $T=57660 48160 0 90 $X=57410 $Y=48080
X86 7 M2_M1_CDNS_9 $T=57670 22770 0 90 $X=57420 $Y=22690
X87 12 M2_M1_CDNS_9 $T=57670 30070 0 90 $X=57420 $Y=29990
X88 6 M2_M1_CDNS_9 $T=57670 37410 0 90 $X=57420 $Y=37330
X89 9 M2_M1_CDNS_9 $T=57670 44710 0 90 $X=57420 $Y=44630
X90 51 M2_M1_CDNS_9 $T=72650 52420 0 90 $X=72400 $Y=52340
X91 35 M2_M1_CDNS_9 $T=78550 36430 0 0 $X=78470 $Y=36180
X92 51 M2_M1_CDNS_9 $T=79400 52420 0 90 $X=79150 $Y=52340
X93 48 M2_M1_CDNS_9 $T=86760 34460 0 0 $X=86680 $Y=34210
X94 49 M2_M1_CDNS_9 $T=86760 49100 0 0 $X=86680 $Y=48850
X95 35 M4_M3_CDNS_12 $T=51080 34160 0 0 $X=51000 $Y=33910
X96 48 M4_M3_CDNS_12 $T=56340 32800 0 0 $X=56260 $Y=32550
X97 49 M4_M3_CDNS_12 $T=56340 47440 0 0 $X=56260 $Y=47190
X98 50 M4_M3_CDNS_12 $T=57240 50840 0 0 $X=57160 $Y=50590
X99 51 M4_M3_CDNS_12 $T=72650 52420 0 90 $X=72400 $Y=52340
X100 35 M4_M3_CDNS_12 $T=78550 36430 0 0 $X=78470 $Y=36180
X101 51 M4_M3_CDNS_12 $T=79400 52420 0 90 $X=79150 $Y=52340
X102 48 M4_M3_CDNS_12 $T=86760 34460 0 0 $X=86680 $Y=34210
X103 49 M4_M3_CDNS_12 $T=86760 49100 0 0 $X=86680 $Y=48850
X104 35 M4_M3_CDNS_13 $T=51140 36930 0 0 $X=51060 $Y=36800
X105 2 M1_PO_CDNS_14 $T=52330 32180 0 90 $X=52080 $Y=32080
X106 35 M1_PO_CDNS_14 $T=52330 46820 0 90 $X=52080 $Y=46720
X107 38 M1_PO_CDNS_14 $T=54270 29810 0 90 $X=54020 $Y=29710
X108 39 M1_PO_CDNS_14 $T=54270 44450 0 90 $X=54020 $Y=44350
X109 36 M1_PO_CDNS_14 $T=55540 26280 0 0 $X=55440 $Y=26030
X110 37 M1_PO_CDNS_14 $T=55540 40920 0 0 $X=55440 $Y=40670
X111 40 M1_PO_CDNS_14 $T=55730 21200 0 90 $X=55480 $Y=21100
X112 41 M1_PO_CDNS_14 $T=55730 35840 0 90 $X=55480 $Y=35740
X113 44 M1_PO_CDNS_14 $T=56050 31070 0 0 $X=55950 $Y=30820
X114 45 M1_PO_CDNS_14 $T=56050 45710 0 0 $X=55950 $Y=45460
X115 42 M1_PO_CDNS_14 $T=56210 23810 0 90 $X=55960 $Y=23710
X116 43 M1_PO_CDNS_14 $T=56210 38450 0 90 $X=55960 $Y=38350
X117 48 M1_PO_CDNS_14 $T=56340 32800 0 0 $X=56240 $Y=32550
X118 49 M1_PO_CDNS_14 $T=56340 47440 0 0 $X=56240 $Y=47190
X119 13 M1_PO_CDNS_14 $T=57660 26200 0 90 $X=57410 $Y=26100
X120 11 M1_PO_CDNS_14 $T=57660 33520 0 90 $X=57410 $Y=33420
X121 10 M1_PO_CDNS_14 $T=57660 40840 0 90 $X=57410 $Y=40740
X122 8 M1_PO_CDNS_14 $T=57660 48160 0 90 $X=57410 $Y=48060
X123 7 M1_PO_CDNS_14 $T=57670 22770 0 90 $X=57420 $Y=22670
X124 12 M1_PO_CDNS_14 $T=57670 30070 0 90 $X=57420 $Y=29970
X125 6 M1_PO_CDNS_14 $T=57670 37410 0 90 $X=57420 $Y=37310
X126 9 M1_PO_CDNS_14 $T=57670 44710 0 90 $X=57420 $Y=44610
X127 35 M1_PO_CDNS_14 $T=78550 36430 0 0 $X=78450 $Y=36180
X128 52 M1_PO_CDNS_15 $T=53520 24980 0 90 $X=53270 $Y=24880
X129 53 M1_PO_CDNS_15 $T=53520 39620 0 90 $X=53270 $Y=39520
X130 14 M1_PO_CDNS_15 $T=64110 23330 0 0 $X=64010 $Y=23080
X131 18 M1_PO_CDNS_15 $T=64110 37970 0 0 $X=64010 $Y=37720
X132 14 M1_PO_CDNS_15 $T=65950 23850 0 90 $X=65700 $Y=23750
X133 18 M1_PO_CDNS_15 $T=65950 38490 0 90 $X=65700 $Y=38390
X134 2 M1_PO_CDNS_15 $T=78510 22370 0 0 $X=78410 $Y=22120
X135 54 M1_PO_CDNS_16 $T=53270 31100 0 0 $X=53170 $Y=30980
X136 55 M1_PO_CDNS_16 $T=53270 45740 0 0 $X=53170 $Y=45620
X137 56 M1_PO_CDNS_16 $T=53550 23450 0 0 $X=53450 $Y=23330
X138 57 M1_PO_CDNS_16 $T=53550 38090 0 0 $X=53450 $Y=37970
X139 58 M1_PO_CDNS_16 $T=53840 25910 0 0 $X=53740 $Y=25790
X140 59 M1_PO_CDNS_16 $T=53840 40550 0 0 $X=53740 $Y=40430
X141 52 M2_M1_CDNS_17 $T=53520 24980 0 90 $X=53270 $Y=24900
X142 53 M2_M1_CDNS_17 $T=53520 39620 0 90 $X=53270 $Y=39540
X143 14 M2_M1_CDNS_17 $T=64110 23330 0 0 $X=64030 $Y=23080
X144 18 M2_M1_CDNS_17 $T=64110 37970 0 0 $X=64030 $Y=37720
X145 14 M2_M1_CDNS_17 $T=65950 23850 0 90 $X=65700 $Y=23770
X146 18 M2_M1_CDNS_17 $T=65950 38490 0 90 $X=65700 $Y=38410
X147 2 M2_M1_CDNS_17 $T=78510 22370 0 0 $X=78430 $Y=22120
X148 3 4 40 56 42 172 NAND_1X_small $T=53960 20720 0 0 $X=53530 $Y=20700
X149 3 4 36 58 52 171 NAND_1X_small $T=55940 28040 0 180 $X=53530 $Y=24260
X150 3 4 38 54 44 170 NAND_1X_small $T=53960 28040 0 0 $X=53530 $Y=28020
X151 3 4 41 57 43 169 NAND_1X_small $T=53960 35360 0 0 $X=53530 $Y=35340
X152 3 4 37 59 53 168 NAND_1X_small $T=55940 42680 0 180 $X=53530 $Y=38900
X153 3 4 39 55 45 167 NAND_1X_small $T=53960 42680 0 0 $X=53530 $Y=42660
X154 3 4 14 7 42 85 86 187 265 188 XOR1 $T=56070 20720 0 0 $X=56130 $Y=20700
X155 3 4 15 13 40 83 84 185 264 186 XOR1 $T=56070 28040 1 0 $X=56130 $Y=24260
X156 3 4 16 12 44 81 82 183 263 184 XOR1 $T=56070 28040 0 0 $X=56130 $Y=28020
X157 3 4 17 11 38 79 80 181 262 182 XOR1 $T=56070 35360 1 0 $X=56130 $Y=31580
X158 3 4 18 6 43 77 78 179 261 180 XOR1 $T=56070 35360 0 0 $X=56130 $Y=35340
X159 3 4 19 10 41 75 76 177 260 178 XOR1 $T=56070 42680 1 0 $X=56130 $Y=38900
X160 3 4 20 9 45 73 74 175 259 176 XOR1 $T=56070 42680 0 0 $X=56130 $Y=42660
X161 3 4 21 8 39 71 72 173 258 174 XOR1 $T=56070 50000 1 0 $X=56130 $Y=46220
X162 5 3 1 4 50 22 51 66 69 70
+ 64 65 67 68 256 257 full_adder1_small $T=50650 49970 0 0 $X=50670 $Y=49980
X163 24 3 23 4 51 33 34 151 154 155
+ 149 150 152 153 266 267 full_adder1_small $T=72610 49970 0 0 $X=72630 $Y=49980
X164 46 48 3 4 2 35 62 63 158 159
+ 254 255 MUX_2to1___2X $T=56190 30160 0 180 $X=50640 $Y=31580
X165 47 49 3 4 35 50 60 61 156 157
+ 252 253 MUX_2to1___2X $T=56190 44800 0 180 $X=50640 $Y=46220
X166 14 13 12 11 3 7 4 15 16 17
+ 2 25 28 27 26 48 140 138 139 FA_4bit $T=64900 20820 0 0 $X=64250 $Y=20700
X167 18 10 9 8 3 6 4 19 20 21
+ 35 32 31 30 29 49 109 107 108 FA_4bit $T=64900 35460 0 0 $X=64250 $Y=35340
X168 56 3 4 52 INV_1X_small $T=51530 20700 0 0 $X=51530 $Y=20700
X169 58 3 4 46 INV_1X_small $T=51530 28060 1 0 $X=51530 $Y=24260
X170 54 3 4 36 INV_1X_small $T=51530 28020 0 0 $X=51530 $Y=28020
X171 57 3 4 53 INV_1X_small $T=51530 35340 0 0 $X=51530 $Y=35340
X172 59 3 4 47 INV_1X_small $T=51530 42700 1 0 $X=51530 $Y=38900
X173 55 3 4 37 INV_1X_small $T=51530 42660 0 0 $X=51530 $Y=42660
M0 64 5 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=16.6612 scb=0.0167915 scc=0.000377457 $X=51440 $Y=52320 $dt=1
M1 58 52 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=25230 $dt=1
M2 59 53 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54550 $Y=39870 $dt=1
M3 56 40 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=23050 $dt=1
M4 54 38 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=30370 $dt=1
M5 57 41 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=37690 $dt=1
M6 55 39 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54850 $Y=45010 $dt=1
M7 3 36 58 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=25230 $dt=1
M8 3 37 59 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=54960 $Y=39870 $dt=1
M9 3 42 56 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=23050 $dt=1
M10 3 44 54 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=30370 $dt=1
M11 3 43 57 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=37690 $dt=1
M12 3 45 55 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=55260 $Y=45010 $dt=1
M13 85 14 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=23040 $dt=1
M14 83 15 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=25240 $dt=1
M15 81 16 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=30360 $dt=1
M16 79 17 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=32560 $dt=1
M17 77 18 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=37680 $dt=1
M18 75 19 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=39880 $dt=1
M19 73 20 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=45000 $dt=1
M20 71 21 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=56900 $Y=47200 $dt=1
M21 86 7 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=23040 $dt=1
M22 84 13 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=25240 $dt=1
M23 82 12 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=30360 $dt=1
M24 80 11 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=32560 $dt=1
M25 78 6 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=37680 $dt=1
M26 76 10 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=39880 $dt=1
M27 74 9 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=45000 $dt=1
M28 72 8 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=57860 $Y=47200 $dt=1
M29 265 7 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=22800 $dt=1
M30 264 13 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=25000 $dt=1
M31 263 12 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=30120 $dt=1
M32 262 11 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=32320 $dt=1
M33 261 6 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=37440 $dt=1
M34 260 10 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=39640 $dt=1
M35 259 9 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=44760 $dt=1
M36 258 8 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=59190 $Y=46960 $dt=1
M37 42 85 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=22860 $dt=1
M38 40 83 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=24940 $dt=1
M39 44 81 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=30180 $dt=1
M40 38 79 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=32260 $dt=1
M41 43 77 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=37500 $dt=1
M42 41 75 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=39580 $dt=1
M43 45 73 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=44820 $dt=1
M44 39 71 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=60160 $Y=46900 $dt=1
M45 42 86 265 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=22860 $dt=1
M46 40 84 264 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=24940 $dt=1
M47 44 82 263 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=30180 $dt=1
M48 38 80 262 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=32260 $dt=1
M49 43 78 261 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=37500 $dt=1
M50 41 76 260 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=39580 $dt=1
M51 45 74 259 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=44820 $dt=1
M52 39 72 258 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.7166 scb=0.00899592 scc=0.000559171 $X=61120 $Y=46900 $dt=1
M53 265 14 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=22860 $dt=1
M54 264 15 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=24940 $dt=1
M55 263 16 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=30180 $dt=1
M56 262 17 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=32260 $dt=1
M57 261 18 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=37500 $dt=1
M58 260 19 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=39580 $dt=1
M59 259 20 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=44820 $dt=1
M60 258 21 3 3 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=15.1061 scb=0.0150932 scc=0.000651875 $X=62080 $Y=46900 $dt=1
M61 34 154 3 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=12.3245 scb=0.0100791 scc=0.000237271 $X=93310 $Y=52330 $dt=1
M62 3 155 34 3 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0172 scb=0.0122201 scc=0.000249942 $X=93720 $Y=52330 $dt=1
.ends 10badder

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_46                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_46 1 2 3 5
*.DEVICECLIMB
** N=5 EP=4 FDC=1
M0 5 3 2 2 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90901 scb=0.00884432 scc=0.000225386 $X=660 $Y=760 $dt=0
.ends cellTmpl_CDNS_46

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: INV_1X_small_layout                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt INV_1X_small_layout 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
X0 1 M1_PO_CDNS_16 $T=700 2040 0 90 $X=580 $Y=1940
X1 2 3 1 4 cellTmpl_CDNS_46 $T=120 140 0 0 $X=0 $Y=0
.ends INV_1X_small_layout

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_clk_part                                  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_clk_part 1 2 3 4 5 6
*.DEVICECLIMB
** N=6 EP=6 FDC=2
X0 1 M1_PO_CDNS_16 $T=640 1830 0 90 $X=520 $Y=1730
X1 6 M1_PO_CDNS_16 $T=1940 640 0 0 $X=1840 $Y=520
X2 3 1 6 3 nmos1v_CDNS_19 $T=710 860 0 0 $X=290 $Y=660
X3 4 6 5 3 nmos1v_CDNS_19 $T=1890 860 0 0 $X=1470 $Y=660
X4 2 3 cellTmpl_CDNS_21 $T=120 140 0 0 $X=0 $Y=0
M0 6 1 3 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=710 $Y=860 $dt=0
M1 5 6 4 3 g45n1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=1890 $Y=860 $dt=0
.ends ph1p3_clk_part

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_48                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_48 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_48

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph1p3_MSDFF                                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph1p3_MSDFF 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17
*.DEVICECLIMB
** N=18 EP=17 FDC=15
X0 7 M3_M2_CDNS_1 $T=1140 2170 0 90 $X=890 $Y=2090
X1 8 M3_M2_CDNS_1 $T=3910 970 0 0 $X=3830 $Y=720
X2 9 M3_M2_CDNS_1 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X3 7 M3_M2_CDNS_1 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X4 7 M3_M2_CDNS_1 $T=8100 2170 0 90 $X=7850 $Y=2090
X5 9 M3_M2_CDNS_1 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X6 8 M3_M2_CDNS_1 $T=9760 1890 0 0 $X=9680 $Y=1640
X7 7 M2_M1_CDNS_2 $T=1140 2170 0 90 $X=890 $Y=2090
X8 8 M2_M1_CDNS_2 $T=3910 970 0 0 $X=3830 $Y=720
X9 9 M2_M1_CDNS_2 $T=4630 -2070 0 0 $X=4550 $Y=-2320
X10 7 M2_M1_CDNS_2 $T=6590 -1760 0 0 $X=6510 $Y=-2010
X11 9 M2_M1_CDNS_2 $T=8890 -1970 0 0 $X=8810 $Y=-2220
X12 8 M2_M1_CDNS_2 $T=9760 1890 0 0 $X=9680 $Y=1640
X13 1 M3_M2_CDNS_7 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X14 1 M3_M2_CDNS_7 $T=5110 3310 0 0 $X=5030 $Y=3060
X15 2 M2_M1_CDNS_8 $T=430 2010 0 0 $X=350 $Y=1880
X16 10 M2_M1_CDNS_8 $T=1110 -1470 0 0 $X=1030 $Y=-1600
X17 2 M2_M1_CDNS_8 $T=2790 -1820 0 0 $X=2710 $Y=-1950
X18 11 M2_M1_CDNS_8 $T=4150 -1460 0 0 $X=4070 $Y=-1590
X19 6 M2_M1_CDNS_8 $T=5200 -2030 0 0 $X=5120 $Y=-2160
X20 10 M2_M1_CDNS_8 $T=5310 1560 0 90 $X=5180 $Y=1480
X21 11 M2_M1_CDNS_8 $T=5670 -1460 0 90 $X=5540 $Y=-1540
X22 12 M2_M1_CDNS_8 $T=6280 1490 0 0 $X=6200 $Y=1360
X23 13 M2_M1_CDNS_8 $T=7300 1510 0 90 $X=7170 $Y=1430
X24 12 M2_M1_CDNS_8 $T=7850 -2080 0 0 $X=7770 $Y=-2210
X25 13 M2_M1_CDNS_8 $T=9400 1510 0 90 $X=9270 $Y=1430
X26 6 M2_M1_CDNS_8 $T=9770 -2060 0 0 $X=9690 $Y=-2190
X27 1 M2_M1_CDNS_9 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X28 1 M2_M1_CDNS_9 $T=5110 3310 0 0 $X=5030 $Y=3060
X29 7 M2_M1_CDNS_9 $T=8100 2170 0 90 $X=7850 $Y=2090
X30 1 M4_M3_CDNS_12 $T=1540 -3270 0 0 $X=1460 $Y=-3520
X31 1 M4_M3_CDNS_12 $T=5110 3310 0 0 $X=5030 $Y=3060
X32 7 M1_PO_CDNS_14 $T=8100 2170 0 90 $X=7850 $Y=2070
X33 8 1 3 10 12 18 NAND2_1X_small $T=3680 -70 0 0 $X=3800 $Y=0
X34 4 1 3 10 INV_1X_small_layout $T=0 40 1 0 $X=0 $Y=-3760
X35 2 1 3 7 INV_1X_small_layout $T=0 0 0 0 $X=0 $Y=0
X36 6 1 3 11 INV_1X_small_layout $T=4800 40 1 0 $X=4800 $Y=-3760
X37 12 1 3 13 INV_1X_small_layout $T=6200 0 0 0 $X=6200 $Y=0
X38 9 1 3 6 INV_1X_small_layout $T=8600 40 1 0 $X=8600 $Y=-3760
X39 2 1 3 5 8 14 ph1p3_clk_part $T=1400 0 0 0 $X=1400 $Y=0
X40 2 1 3 11 9 15 ph1p3_clk_part $T=2400 40 1 0 $X=2400 $Y=-3760
X41 7 1 3 12 9 16 ph1p3_clk_part $T=6200 40 1 0 $X=6200 $Y=-3760
X42 7 1 3 13 8 17 ph1p3_clk_part $T=7600 0 0 0 $X=7600 $Y=0
X43 1 3 cellTmpl_CDNS_48 $T=1520 -100 1 0 $X=1400 $Y=-3760
.ends ph1p3_MSDFF

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: cellTmpl_CDNS_49                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt cellTmpl_CDNS_49 1 2
** N=2 EP=2 FDC=0
.ends cellTmpl_CDNS_49

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MUX_2to1___2X_ph2p2                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MUX_2to1___2X_ph2p2 1 2 3 4 5 6 7 8 9 10
+ 11 12
*.DEVICECLIMB
** N=12 EP=12 FDC=6
X0 7 M3_M2_CDNS_1 $T=430 2220 0 0 $X=350 $Y=1970
X1 7 M3_M2_CDNS_1 $T=1140 3180 0 0 $X=1060 $Y=2930
X2 7 M3_M2_CDNS_1 $T=2800 2490 0 0 $X=2720 $Y=2240
X3 7 M2_M1_CDNS_2 $T=1140 3180 0 0 $X=1060 $Y=2930
X4 7 M2_M1_CDNS_9 $T=430 2220 0 0 $X=350 $Y=1970
X5 7 M2_M1_CDNS_9 $T=2800 2490 0 0 $X=2720 $Y=2240
X6 7 M1_PO_CDNS_14 $T=430 2220 0 0 $X=330 $Y=1970
X7 7 M1_PO_CDNS_14 $T=2800 2490 0 0 $X=2700 $Y=2240
X8 1 M1_PO_CDNS_15 $T=1480 1720 0 0 $X=1380 $Y=1470
X9 1 M1_PO_CDNS_15 $T=2840 980 0 0 $X=2740 $Y=730
X10 1 M1_PO_CDNS_16 $T=860 1670 0 0 $X=760 $Y=1550
X11 2 M1_PO_CDNS_16 $T=1480 3130 0 0 $X=1380 $Y=3010
X12 5 M1_PO_CDNS_16 $T=4220 2040 0 0 $X=4120 $Y=1920
X13 8 M1_PO_CDNS_16 $T=4480 1550 0 90 $X=4360 $Y=1450
X14 1 M2_M1_CDNS_17 $T=1480 1720 0 0 $X=1400 $Y=1470
X15 1 M2_M1_CDNS_17 $T=2840 980 0 0 $X=2760 $Y=730
X16 4 7 9 4 nmos1v_CDNS_31 $T=2170 800 0 0 $X=1970 $Y=600
X17 8 5 10 4 nmos1v_CDNS_31 $T=3550 790 0 0 $X=3350 $Y=590
X18 8 2 9 4 nmos1v_CDNS_32 $T=1960 800 0 0 $X=1540 $Y=600
X19 4 1 10 4 nmos1v_CDNS_32 $T=3340 790 0 0 $X=2920 $Y=590
X20 3 4 1 7 8 6 cellTmpl_CDNS_43 $T=120 140 0 0 $X=0 $Y=0
X21 3 1 11 4 3 pmos1v_CDNS_44 $T=2170 2100 0 0 $X=1970 $Y=1900
X22 8 5 12 4 3 pmos1v_CDNS_44 $T=3550 2030 0 0 $X=3350 $Y=1830
X23 8 2 11 4 3 pmos1v_CDNS_45 $T=1960 2100 0 0 $X=1540 $Y=1900
X24 3 7 12 4 3 pmos1v_CDNS_45 $T=3340 2030 0 0 $X=2920 $Y=1830
M0 9 2 8 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=1960 $Y=800 $dt=0
M1 4 7 9 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.8836 scb=0.0102333 scc=0.000414887 $X=2170 $Y=800 $dt=0
M2 10 1 4 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=1.44e-14 AS=3.36e-14 PD=6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=2.45e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3340 $Y=790 $dt=0
M3 8 5 10 4 g45n1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=1.44e-14 PD=7.6e-07 PS=6e-07 fw=2.4e-07 sa=2.45e-07 sb=1.4e-07 sca=10.6427 scb=0.00988663 scc=0.000381704 $X=3550 $Y=790 $dt=0
.ends MUX_2to1___2X_ph2p2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p2_processing_element                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p2_processing_element 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 77 78 79 81 83
+ 108 113 130 139 140 141 158 159 176 185
+ 190 191 194 211 212 213 330 332 333 334
+ 336 338 348 350 351 352 354 356 366 368
+ 369 370 372 374 505 691 697 703 760 761
+ 762 763
*.DEVICECLIMB
** N=789 EP=122 FDC=1597
X0 6 M3_M2_CDNS_1 $T=1860 60810 0 0 $X=1780 $Y=60560
X1 6 M3_M2_CDNS_1 $T=1870 68120 0 0 $X=1790 $Y=67870
X2 6 M3_M2_CDNS_1 $T=12100 60800 0 0 $X=12020 $Y=60550
X3 6 M3_M2_CDNS_1 $T=12100 68120 0 0 $X=12020 $Y=67870
X4 6 M3_M2_CDNS_1 $T=22340 68120 0 0 $X=22260 $Y=67870
X5 6 M3_M2_CDNS_1 $T=22350 60800 0 0 $X=22270 $Y=60550
X6 46 M3_M2_CDNS_1 $T=22980 34240 0 0 $X=22900 $Y=33990
X7 47 M3_M2_CDNS_1 $T=28400 24370 0 0 $X=28320 $Y=24120
X8 48 M3_M2_CDNS_1 $T=32190 56290 0 0 $X=32110 $Y=56040
X9 6 M3_M2_CDNS_1 $T=32580 60800 0 0 $X=32500 $Y=60550
X10 6 M3_M2_CDNS_1 $T=32580 68120 0 0 $X=32500 $Y=67870
X11 6 M3_M2_CDNS_1 $T=40360 10220 0 90 $X=40110 $Y=10140
X12 6 M3_M2_CDNS_1 $T=40340 24940 0 0 $X=40260 $Y=24690
X13 6 M3_M2_CDNS_1 $T=40370 17590 0 0 $X=40290 $Y=17340
X14 49 M3_M2_CDNS_1 $T=45710 34580 0 0 $X=45630 $Y=34330
X15 6 M3_M2_CDNS_1 $T=47620 54480 0 90 $X=47370 $Y=54400
X16 6 M3_M2_CDNS_1 $T=47800 38230 0 90 $X=47550 $Y=38150
X17 6 M3_M2_CDNS_1 $T=47870 10240 0 0 $X=47790 $Y=9990
X18 6 M3_M2_CDNS_1 $T=48260 51950 0 90 $X=48010 $Y=51870
X19 6 M3_M2_CDNS_1 $T=48260 45130 0 0 $X=48180 $Y=44880
X20 6 M3_M2_CDNS_1 $T=48690 16910 0 0 $X=48610 $Y=16660
X21 6 M3_M2_CDNS_1 $T=48860 24230 0 0 $X=48780 $Y=23980
X22 50 M2_M1_CDNS_2 $T=14700 34240 0 0 $X=14620 $Y=33990
X23 46 M2_M1_CDNS_2 $T=22980 34240 0 0 $X=22900 $Y=33990
X24 47 M2_M1_CDNS_2 $T=28400 24370 0 0 $X=28320 $Y=24120
X25 48 M2_M1_CDNS_2 $T=32190 56290 0 0 $X=32110 $Y=56040
X26 51 M2_M1_CDNS_2 $T=38820 45300 0 0 $X=38740 $Y=45050
X27 49 M2_M1_CDNS_2 $T=45710 34580 0 0 $X=45630 $Y=34330
X28 52 M4_M3_CDNS_3 $T=32380 35710 0 90 $X=32130 $Y=35630
X29 53 M4_M3_CDNS_3 $T=33360 32510 0 90 $X=33110 $Y=32430
X30 54 M4_M3_CDNS_3 $T=33880 28620 0 0 $X=33800 $Y=28370
X31 55 M4_M3_CDNS_3 $T=34010 30140 0 0 $X=33930 $Y=29890
X32 56 M4_M3_CDNS_3 $T=34370 21060 0 0 $X=34290 $Y=20810
X33 57 M4_M3_CDNS_3 $T=36160 20250 0 0 $X=36080 $Y=20000
X34 58 M4_M3_CDNS_3 $T=36500 13950 0 0 $X=36420 $Y=13700
X35 59 M4_M3_CDNS_3 $T=37400 32460 0 0 $X=37320 $Y=32210
X36 60 M4_M3_CDNS_3 $T=37820 20120 0 0 $X=37740 $Y=19870
X37 58 M4_M3_CDNS_3 $T=40460 17040 0 90 $X=40210 $Y=16960
X38 60 M4_M3_CDNS_3 $T=40660 20120 0 90 $X=40410 $Y=20040
X39 61 M4_M3_CDNS_3 $T=40730 9730 0 90 $X=40480 $Y=9650
X40 62 M4_M3_CDNS_3 $T=40560 26320 0 0 $X=40480 $Y=26070
X41 59 M4_M3_CDNS_3 $T=42630 35130 0 90 $X=42380 $Y=35050
X42 7 M4_M3_CDNS_3 $T=47890 45870 0 0 $X=47810 $Y=45620
X43 63 M3_M2_CDNS_4 $T=14040 560 0 0 $X=13960 $Y=430
X44 64 M3_M2_CDNS_4 $T=22250 3160 0 0 $X=22170 $Y=3030
X45 63 M3_M2_CDNS_4 $T=23920 6540 0 0 $X=23840 $Y=6410
X46 48 M3_M2_CDNS_4 $T=25520 48970 0 0 $X=25440 $Y=48840
X47 65 M3_M2_CDNS_4 $T=27740 16660 0 0 $X=27660 $Y=16530
X48 51 M3_M2_CDNS_4 $T=28010 24010 0 0 $X=27930 $Y=23880
X49 59 M3_M2_CDNS_4 $T=31460 30680 0 90 $X=31330 $Y=30600
X50 48 M3_M2_CDNS_4 $T=32190 54030 0 0 $X=32110 $Y=53900
X51 53 M3_M2_CDNS_4 $T=36910 32510 0 0 $X=36830 $Y=32380
X52 53 M3_M2_CDNS_4 $T=37470 13030 0 0 $X=37390 $Y=12900
X53 66 M3_M2_CDNS_4 $T=37590 8380 0 90 $X=37460 $Y=8300
X54 66 M3_M2_CDNS_4 $T=38080 28430 0 0 $X=38000 $Y=28300
X55 49 M3_M2_CDNS_4 $T=39590 33870 0 0 $X=39510 $Y=33740
X56 52 M3_M2_CDNS_4 $T=40110 35670 0 90 $X=39980 $Y=35590
X57 67 M3_M2_CDNS_4 $T=42020 34330 0 0 $X=41940 $Y=34200
X58 54 M3_M2_CDNS_4 $T=45640 37660 0 0 $X=45560 $Y=37530
X59 6 M3_M2_CDNS_4 $T=47780 30450 0 0 $X=47700 $Y=30320
X60 6 M3_M2_CDNS_4 $T=47810 35930 0 0 $X=47730 $Y=35800
X61 60 M3_M2_CDNS_4 $T=48170 20860 0 0 $X=48090 $Y=20730
X62 62 M3_M2_CDNS_4 $T=48180 28260 0 0 $X=48100 $Y=28130
X63 7 M3_M2_CDNS_4 $T=48350 54060 0 0 $X=48270 $Y=53930
X64 58 M3_M2_CDNS_4 $T=48430 15830 0 0 $X=48350 $Y=15700
X65 59 M3_M2_CDNS_4 $T=49580 57720 0 90 $X=49450 $Y=57640
X66 61 M3_M2_CDNS_4 $T=50600 8490 0 0 $X=50520 $Y=8360
X67 1 M5_M4_CDNS_5 $T=1480 56760 0 0 $X=1400 $Y=56510
X68 4 M5_M4_CDNS_5 $T=2350 44590 0 90 $X=2100 $Y=44510
X69 3 M5_M4_CDNS_5 $T=3900 48300 0 90 $X=3650 $Y=48220
X70 2 M5_M4_CDNS_5 $T=3940 58210 0 90 $X=3690 $Y=58130
X71 1 M5_M4_CDNS_5 $T=4250 65060 0 0 $X=4170 $Y=64810
X72 2 M5_M4_CDNS_5 $T=4250 72470 0 0 $X=4170 $Y=72220
X73 11 M5_M4_CDNS_5 $T=6840 58120 0 90 $X=6590 $Y=58040
X74 15 M5_M4_CDNS_5 $T=11380 56560 0 90 $X=11130 $Y=56480
X75 15 M5_M4_CDNS_5 $T=14490 65150 0 0 $X=14410 $Y=64900
X76 11 M5_M4_CDNS_5 $T=14490 72480 0 0 $X=14410 $Y=72230
X77 14 M5_M4_CDNS_5 $T=20420 56560 0 90 $X=20170 $Y=56480
X78 14 M5_M4_CDNS_5 $T=24730 65150 0 0 $X=24650 $Y=64900
X79 3 M5_M4_CDNS_5 $T=24730 72470 0 0 $X=24650 $Y=72220
X80 52 M5_M4_CDNS_5 $T=27620 26990 0 0 $X=27540 $Y=26740
X81 16 M5_M4_CDNS_5 $T=29230 56560 0 90 $X=28980 $Y=56480
X82 52 M5_M4_CDNS_5 $T=32380 35710 0 90 $X=32130 $Y=35630
X83 53 M5_M4_CDNS_5 $T=32470 34080 0 90 $X=32220 $Y=34000
X84 53 M5_M4_CDNS_5 $T=33360 32510 0 90 $X=33110 $Y=32430
X85 68 M5_M4_CDNS_5 $T=33670 6150 0 90 $X=33420 $Y=6070
X86 54 M5_M4_CDNS_5 $T=33880 28620 0 0 $X=33800 $Y=28370
X87 55 M5_M4_CDNS_5 $T=34010 30140 0 0 $X=33930 $Y=29890
X88 56 M5_M4_CDNS_5 $T=34370 21060 0 0 $X=34290 $Y=20810
X89 16 M5_M4_CDNS_5 $T=34970 65150 0 0 $X=34890 $Y=64900
X90 4 M5_M4_CDNS_5 $T=34970 72470 0 0 $X=34890 $Y=72220
X91 55 M5_M4_CDNS_5 $T=35130 53970 0 0 $X=35050 $Y=53720
X92 57 M5_M4_CDNS_5 $T=36160 20250 0 0 $X=36080 $Y=20000
X93 58 M5_M4_CDNS_5 $T=36500 13950 0 0 $X=36420 $Y=13700
X94 59 M5_M4_CDNS_5 $T=37400 32460 0 0 $X=37320 $Y=32210
X95 60 M5_M4_CDNS_5 $T=37820 20120 0 0 $X=37740 $Y=19870
X96 63 M5_M4_CDNS_5 $T=38220 15840 0 0 $X=38140 $Y=15590
X97 68 M5_M4_CDNS_5 $T=38250 22590 0 0 $X=38170 $Y=22340
X98 57 M5_M4_CDNS_5 $T=38270 21170 0 0 $X=38190 $Y=20920
X99 58 M5_M4_CDNS_5 $T=40460 17040 0 90 $X=40210 $Y=16960
X100 60 M5_M4_CDNS_5 $T=40660 20120 0 90 $X=40410 $Y=20040
X101 61 M5_M4_CDNS_5 $T=40730 9730 0 90 $X=40480 $Y=9650
X102 62 M5_M4_CDNS_5 $T=40560 26320 0 0 $X=40480 $Y=26070
X103 59 M5_M4_CDNS_5 $T=42630 35130 0 90 $X=42380 $Y=35050
X104 69 M5_M4_CDNS_5 $T=47280 7640 0 90 $X=47030 $Y=7560
X105 63 M5_M4_CDNS_5 $T=47850 15290 0 0 $X=47770 $Y=15040
X106 68 M5_M4_CDNS_5 $T=47850 23870 0 0 $X=47770 $Y=23620
X107 7 M5_M4_CDNS_5 $T=47890 45870 0 0 $X=47810 $Y=45620
X108 6 M5_M4_CDNS_5 $T=47980 9490 0 0 $X=47900 $Y=9240
X109 6 M5_M4_CDNS_5 $T=48880 2280 0 0 $X=48800 $Y=2030
X110 7 M5_M4_CDNS_5 $T=50250 45640 0 90 $X=50000 $Y=45560
X111 69 M5_M4_CDNS_5 $T=59660 13790 0 0 $X=59580 $Y=13540
X112 63 M5_M4_CDNS_5 $T=59660 21120 0 0 $X=59580 $Y=20870
X113 68 M5_M4_CDNS_5 $T=59660 28470 0 0 $X=59580 $Y=28220
X114 1 M4_M3_CDNS_6 $T=1480 56760 0 0 $X=1400 $Y=56510
X115 4 M4_M3_CDNS_6 $T=2350 44590 0 90 $X=2100 $Y=44510
X116 3 M4_M3_CDNS_6 $T=3900 48300 0 90 $X=3650 $Y=48220
X117 2 M4_M3_CDNS_6 $T=3940 58210 0 90 $X=3690 $Y=58130
X118 1 M4_M3_CDNS_6 $T=4250 65060 0 0 $X=4170 $Y=64810
X119 2 M4_M3_CDNS_6 $T=4250 72470 0 0 $X=4170 $Y=72220
X120 11 M4_M3_CDNS_6 $T=6840 58120 0 90 $X=6590 $Y=58040
X121 15 M4_M3_CDNS_6 $T=11380 56560 0 90 $X=11130 $Y=56480
X122 15 M4_M3_CDNS_6 $T=14490 65150 0 0 $X=14410 $Y=64900
X123 11 M4_M3_CDNS_6 $T=14490 72480 0 0 $X=14410 $Y=72230
X124 14 M4_M3_CDNS_6 $T=20420 56560 0 90 $X=20170 $Y=56480
X125 14 M4_M3_CDNS_6 $T=24730 65150 0 0 $X=24650 $Y=64900
X126 3 M4_M3_CDNS_6 $T=24730 72470 0 0 $X=24650 $Y=72220
X127 52 M4_M3_CDNS_6 $T=27620 26990 0 0 $X=27540 $Y=26740
X128 16 M4_M3_CDNS_6 $T=29230 56560 0 90 $X=28980 $Y=56480
X129 53 M4_M3_CDNS_6 $T=32470 34080 0 90 $X=32220 $Y=34000
X130 68 M4_M3_CDNS_6 $T=33670 6150 0 90 $X=33420 $Y=6070
X131 16 M4_M3_CDNS_6 $T=34970 65150 0 0 $X=34890 $Y=64900
X132 4 M4_M3_CDNS_6 $T=34970 72470 0 0 $X=34890 $Y=72220
X133 55 M4_M3_CDNS_6 $T=35130 53970 0 0 $X=35050 $Y=53720
X134 63 M4_M3_CDNS_6 $T=38220 15840 0 0 $X=38140 $Y=15590
X135 68 M4_M3_CDNS_6 $T=38250 22590 0 0 $X=38170 $Y=22340
X136 57 M4_M3_CDNS_6 $T=38270 21170 0 0 $X=38190 $Y=20920
X137 69 M4_M3_CDNS_6 $T=47280 7640 0 90 $X=47030 $Y=7560
X138 63 M4_M3_CDNS_6 $T=47850 15290 0 0 $X=47770 $Y=15040
X139 68 M4_M3_CDNS_6 $T=47850 23870 0 0 $X=47770 $Y=23620
X140 6 M4_M3_CDNS_6 $T=47980 9490 0 0 $X=47900 $Y=9240
X141 6 M4_M3_CDNS_6 $T=48880 2280 0 0 $X=48800 $Y=2030
X142 7 M4_M3_CDNS_6 $T=50250 45640 0 90 $X=50000 $Y=45560
X143 69 M4_M3_CDNS_6 $T=59660 13790 0 0 $X=59580 $Y=13540
X144 63 M4_M3_CDNS_6 $T=59660 21120 0 0 $X=59580 $Y=20870
X145 68 M4_M3_CDNS_6 $T=59660 28470 0 0 $X=59580 $Y=28220
X146 5 M3_M2_CDNS_7 $T=1340 55390 0 0 $X=1260 $Y=55140
X147 1 M3_M2_CDNS_7 $T=1480 56760 0 0 $X=1400 $Y=56510
X148 4 M3_M2_CDNS_7 $T=2350 44590 0 90 $X=2100 $Y=44510
X149 5 M3_M2_CDNS_7 $T=3450 61970 0 0 $X=3370 $Y=61720
X150 3 M3_M2_CDNS_7 $T=3900 48300 0 90 $X=3650 $Y=48220
X151 2 M3_M2_CDNS_7 $T=3940 58210 0 90 $X=3690 $Y=58130
X152 1 M3_M2_CDNS_7 $T=4250 65060 0 0 $X=4170 $Y=64810
X153 2 M3_M2_CDNS_7 $T=4250 72470 0 0 $X=4170 $Y=72220
X154 11 M3_M2_CDNS_7 $T=6840 58120 0 90 $X=6590 $Y=58040
X155 5 M3_M2_CDNS_7 $T=9870 69280 0 0 $X=9790 $Y=69030
X156 15 M3_M2_CDNS_7 $T=11380 56560 0 90 $X=11130 $Y=56480
X157 15 M3_M2_CDNS_7 $T=14490 65150 0 0 $X=14410 $Y=64900
X158 11 M3_M2_CDNS_7 $T=14490 72480 0 0 $X=14410 $Y=72230
X159 50 M3_M2_CDNS_7 $T=14700 34240 0 0 $X=14620 $Y=33990
X160 14 M3_M2_CDNS_7 $T=20420 56560 0 90 $X=20170 $Y=56480
X161 14 M3_M2_CDNS_7 $T=24730 65150 0 0 $X=24650 $Y=64900
X162 3 M3_M2_CDNS_7 $T=24730 72470 0 0 $X=24650 $Y=72220
X163 52 M3_M2_CDNS_7 $T=27620 26990 0 0 $X=27540 $Y=26740
X164 67 M3_M2_CDNS_7 $T=28040 20980 0 0 $X=27960 $Y=20730
X165 16 M3_M2_CDNS_7 $T=29230 56560 0 90 $X=28980 $Y=56480
X166 53 M3_M2_CDNS_7 $T=32470 34080 0 90 $X=32220 $Y=34000
X167 68 M3_M2_CDNS_7 $T=33670 6150 0 90 $X=33420 $Y=6070
X168 16 M3_M2_CDNS_7 $T=34970 65150 0 0 $X=34890 $Y=64900
X169 4 M3_M2_CDNS_7 $T=34970 72470 0 0 $X=34890 $Y=72220
X170 55 M3_M2_CDNS_7 $T=35130 53970 0 0 $X=35050 $Y=53720
X171 49 M3_M2_CDNS_7 $T=37620 30320 0 0 $X=37540 $Y=30070
X172 63 M3_M2_CDNS_7 $T=38220 15840 0 0 $X=38140 $Y=15590
X173 68 M3_M2_CDNS_7 $T=38250 22590 0 0 $X=38170 $Y=22340
X174 57 M3_M2_CDNS_7 $T=38270 21170 0 0 $X=38190 $Y=20920
X175 51 M3_M2_CDNS_7 $T=38820 45300 0 0 $X=38740 $Y=45050
X176 70 M3_M2_CDNS_7 $T=40600 13810 0 0 $X=40520 $Y=13560
X177 64 M3_M2_CDNS_7 $T=40710 21060 0 0 $X=40630 $Y=20810
X178 7 M3_M2_CDNS_7 $T=46890 13630 0 0 $X=46810 $Y=13380
X179 7 M3_M2_CDNS_7 $T=46900 20740 0 0 $X=46820 $Y=20490
X180 7 M3_M2_CDNS_7 $T=46910 28080 0 0 $X=46830 $Y=27830
X181 69 M3_M2_CDNS_7 $T=47280 7640 0 90 $X=47030 $Y=7560
X182 63 M3_M2_CDNS_7 $T=47850 15290 0 0 $X=47770 $Y=15040
X183 68 M3_M2_CDNS_7 $T=47850 23870 0 0 $X=47770 $Y=23620
X184 6 M3_M2_CDNS_7 $T=47980 9490 0 0 $X=47900 $Y=9240
X185 6 M3_M2_CDNS_7 $T=48880 2280 0 0 $X=48800 $Y=2030
X186 5 M3_M2_CDNS_7 $T=49180 4060 0 0 $X=49100 $Y=3810
X187 5 M3_M2_CDNS_7 $T=49180 11470 0 0 $X=49100 $Y=11220
X188 5 M3_M2_CDNS_7 $T=49180 18800 0 0 $X=49100 $Y=18550
X189 5 M3_M2_CDNS_7 $T=49180 26120 0 0 $X=49100 $Y=25870
X190 5 M3_M2_CDNS_7 $T=49180 33430 0 0 $X=49100 $Y=33180
X191 5 M3_M2_CDNS_7 $T=49180 40820 0 0 $X=49100 $Y=40570
X192 5 M3_M2_CDNS_7 $T=49180 48070 0 0 $X=49100 $Y=47820
X193 5 M3_M2_CDNS_7 $T=49180 54710 0 0 $X=49100 $Y=54460
X194 7 M3_M2_CDNS_7 $T=50250 45640 0 90 $X=50000 $Y=45560
X195 71 M3_M2_CDNS_7 $T=50910 13780 0 0 $X=50830 $Y=13530
X196 25 M3_M2_CDNS_7 $T=58670 9650 0 90 $X=58420 $Y=9570
X197 25 M3_M2_CDNS_7 $T=58670 12550 0 90 $X=58420 $Y=12470
X198 25 M3_M2_CDNS_7 $T=58670 16970 0 90 $X=58420 $Y=16890
X199 25 M3_M2_CDNS_7 $T=58670 19870 0 90 $X=58420 $Y=19790
X200 25 M3_M2_CDNS_7 $T=58670 24290 0 90 $X=58420 $Y=24210
X201 25 M3_M2_CDNS_7 $T=58670 27190 0 90 $X=58420 $Y=27110
X202 25 M3_M2_CDNS_7 $T=58670 31610 0 90 $X=58420 $Y=31530
X203 25 M3_M2_CDNS_7 $T=58670 38930 0 90 $X=58420 $Y=38850
X204 25 M3_M2_CDNS_7 $T=58670 46250 0 90 $X=58420 $Y=46170
X205 25 M3_M2_CDNS_7 $T=58670 53570 0 90 $X=58420 $Y=53490
X206 69 M3_M2_CDNS_7 $T=59660 13790 0 0 $X=59580 $Y=13540
X207 63 M3_M2_CDNS_7 $T=59660 21120 0 0 $X=59580 $Y=20870
X208 68 M3_M2_CDNS_7 $T=59660 28470 0 0 $X=59580 $Y=28220
X209 64 M2_M1_CDNS_8 $T=13960 1790 0 90 $X=13830 $Y=1710
X210 72 M2_M1_CDNS_8 $T=26670 45180 0 0 $X=26590 $Y=45050
X211 59 M2_M1_CDNS_8 $T=27600 31220 0 0 $X=27520 $Y=31090
X212 66 M2_M1_CDNS_8 $T=28050 6240 0 0 $X=27970 $Y=6110
X213 60 M2_M1_CDNS_8 $T=28100 13310 0 0 $X=28020 $Y=13180
X214 71 M2_M1_CDNS_8 $T=28110 10050 0 0 $X=28030 $Y=9920
X215 62 M2_M1_CDNS_8 $T=28410 16430 0 90 $X=28280 $Y=16350
X216 53 M2_M1_CDNS_8 $T=35470 34490 0 0 $X=35390 $Y=34360
X217 70 M2_M1_CDNS_8 $T=35820 2210 0 90 $X=35690 $Y=2130
X218 65 M2_M1_CDNS_8 $T=37240 38080 0 0 $X=37160 $Y=37950
X219 66 M2_M1_CDNS_8 $T=41060 27730 0 0 $X=40980 $Y=27600
X220 73 M2_M1_CDNS_8 $T=43080 53380 0 0 $X=43000 $Y=53250
X221 7 M2_M1_CDNS_8 $T=47420 36740 0 0 $X=47340 $Y=36610
X222 49 M2_M1_CDNS_8 $T=47770 37090 0 0 $X=47690 $Y=36960
X223 52 M2_M1_CDNS_8 $T=50960 49840 0 90 $X=50830 $Y=49760
X224 47 M2_M1_CDNS_8 $T=51290 41540 0 90 $X=51160 $Y=41460
X225 60 M2_M1_CDNS_8 $T=51280 20630 0 0 $X=51200 $Y=20500
X226 67 M2_M1_CDNS_8 $T=51290 35200 0 0 $X=51210 $Y=35070
X227 62 M2_M1_CDNS_8 $T=51300 27960 0 0 $X=51220 $Y=27830
X228 59 M2_M1_CDNS_8 $T=51300 57100 0 0 $X=51220 $Y=56970
X229 61 M2_M1_CDNS_8 $T=59660 8330 0 0 $X=59580 $Y=8200
X230 58 M2_M1_CDNS_8 $T=59660 15640 0 0 $X=59580 $Y=15510
X231 57 M2_M1_CDNS_8 $T=59660 22940 0 0 $X=59580 $Y=22810
X232 56 M2_M1_CDNS_8 $T=59660 30310 0 0 $X=59580 $Y=30180
X233 49 M2_M1_CDNS_8 $T=59660 37620 0 0 $X=59580 $Y=37490
X234 54 M2_M1_CDNS_8 $T=59660 44940 0 0 $X=59580 $Y=44810
X235 55 M2_M1_CDNS_8 $T=59660 52270 0 0 $X=59580 $Y=52140
X236 5 M2_M1_CDNS_9 $T=1340 55390 0 0 $X=1260 $Y=55140
X237 1 M2_M1_CDNS_9 $T=1480 56760 0 0 $X=1400 $Y=56510
X238 6 M2_M1_CDNS_9 $T=1860 60810 0 0 $X=1780 $Y=60560
X239 6 M2_M1_CDNS_9 $T=1870 68120 0 0 $X=1790 $Y=67870
X240 4 M2_M1_CDNS_9 $T=2350 44590 0 90 $X=2100 $Y=44510
X241 5 M2_M1_CDNS_9 $T=3450 61970 0 0 $X=3370 $Y=61720
X242 3 M2_M1_CDNS_9 $T=3900 48300 0 90 $X=3650 $Y=48220
X243 2 M2_M1_CDNS_9 $T=3940 58210 0 90 $X=3690 $Y=58130
X244 1 M2_M1_CDNS_9 $T=4250 65060 0 0 $X=4170 $Y=64810
X245 2 M2_M1_CDNS_9 $T=4250 72470 0 0 $X=4170 $Y=72220
X246 11 M2_M1_CDNS_9 $T=6840 58120 0 90 $X=6590 $Y=58040
X247 5 M2_M1_CDNS_9 $T=9870 69280 0 0 $X=9790 $Y=69030
X248 15 M2_M1_CDNS_9 $T=11380 56560 0 90 $X=11130 $Y=56480
X249 6 M2_M1_CDNS_9 $T=12100 60800 0 0 $X=12020 $Y=60550
X250 6 M2_M1_CDNS_9 $T=12100 68120 0 0 $X=12020 $Y=67870
X251 15 M2_M1_CDNS_9 $T=14490 65150 0 0 $X=14410 $Y=64900
X252 11 M2_M1_CDNS_9 $T=14490 72480 0 0 $X=14410 $Y=72230
X253 14 M2_M1_CDNS_9 $T=20420 56560 0 90 $X=20170 $Y=56480
X254 6 M2_M1_CDNS_9 $T=22340 68120 0 0 $X=22260 $Y=67870
X255 6 M2_M1_CDNS_9 $T=22350 60800 0 0 $X=22270 $Y=60550
X256 14 M2_M1_CDNS_9 $T=24730 65150 0 0 $X=24650 $Y=64900
X257 3 M2_M1_CDNS_9 $T=24730 72470 0 0 $X=24650 $Y=72220
X258 52 M2_M1_CDNS_9 $T=27620 26990 0 0 $X=27540 $Y=26740
X259 67 M2_M1_CDNS_9 $T=28040 20980 0 0 $X=27960 $Y=20730
X260 16 M2_M1_CDNS_9 $T=29230 56560 0 90 $X=28980 $Y=56480
X261 6 M2_M1_CDNS_9 $T=32580 60800 0 0 $X=32500 $Y=60550
X262 6 M2_M1_CDNS_9 $T=32580 68120 0 0 $X=32500 $Y=67870
X263 68 M2_M1_CDNS_9 $T=33670 6150 0 90 $X=33420 $Y=6070
X264 16 M2_M1_CDNS_9 $T=34970 65150 0 0 $X=34890 $Y=64900
X265 4 M2_M1_CDNS_9 $T=34970 72470 0 0 $X=34890 $Y=72220
X266 49 M2_M1_CDNS_9 $T=37620 30320 0 0 $X=37540 $Y=30070
X267 6 M2_M1_CDNS_9 $T=40360 10220 0 90 $X=40110 $Y=10140
X268 6 M2_M1_CDNS_9 $T=40340 24940 0 0 $X=40260 $Y=24690
X269 6 M2_M1_CDNS_9 $T=40370 17590 0 0 $X=40290 $Y=17340
X270 70 M2_M1_CDNS_9 $T=40600 13810 0 0 $X=40520 $Y=13560
X271 64 M2_M1_CDNS_9 $T=40710 21060 0 0 $X=40630 $Y=20810
X272 7 M2_M1_CDNS_9 $T=46890 13630 0 0 $X=46810 $Y=13380
X273 7 M2_M1_CDNS_9 $T=46900 20740 0 0 $X=46820 $Y=20490
X274 7 M2_M1_CDNS_9 $T=46910 28080 0 0 $X=46830 $Y=27830
X275 6 M2_M1_CDNS_9 $T=47620 54480 0 90 $X=47370 $Y=54400
X276 6 M2_M1_CDNS_9 $T=47800 38230 0 90 $X=47550 $Y=38150
X277 6 M2_M1_CDNS_9 $T=47870 10240 0 0 $X=47790 $Y=9990
X278 6 M2_M1_CDNS_9 $T=47980 9490 0 0 $X=47900 $Y=9240
X279 6 M2_M1_CDNS_9 $T=48260 51950 0 90 $X=48010 $Y=51870
X280 6 M2_M1_CDNS_9 $T=48260 45130 0 0 $X=48180 $Y=44880
X281 6 M2_M1_CDNS_9 $T=48690 16910 0 0 $X=48610 $Y=16660
X282 6 M2_M1_CDNS_9 $T=48860 24230 0 0 $X=48780 $Y=23980
X283 6 M2_M1_CDNS_9 $T=48880 2280 0 0 $X=48800 $Y=2030
X284 5 M2_M1_CDNS_9 $T=49180 4060 0 0 $X=49100 $Y=3810
X285 5 M2_M1_CDNS_9 $T=49180 11470 0 0 $X=49100 $Y=11220
X286 5 M2_M1_CDNS_9 $T=49180 18800 0 0 $X=49100 $Y=18550
X287 5 M2_M1_CDNS_9 $T=49180 26120 0 0 $X=49100 $Y=25870
X288 5 M2_M1_CDNS_9 $T=49180 33430 0 0 $X=49100 $Y=33180
X289 5 M2_M1_CDNS_9 $T=49180 40820 0 0 $X=49100 $Y=40570
X290 5 M2_M1_CDNS_9 $T=49180 48070 0 0 $X=49100 $Y=47820
X291 5 M2_M1_CDNS_9 $T=49180 54710 0 0 $X=49100 $Y=54460
X292 71 M2_M1_CDNS_9 $T=50910 13780 0 0 $X=50830 $Y=13530
X293 25 M2_M1_CDNS_9 $T=58670 9650 0 90 $X=58420 $Y=9570
X294 25 M2_M1_CDNS_9 $T=58670 12550 0 90 $X=58420 $Y=12470
X295 25 M2_M1_CDNS_9 $T=58670 16970 0 90 $X=58420 $Y=16890
X296 25 M2_M1_CDNS_9 $T=58670 19870 0 90 $X=58420 $Y=19790
X297 25 M2_M1_CDNS_9 $T=58670 24290 0 90 $X=58420 $Y=24210
X298 25 M2_M1_CDNS_9 $T=58670 27190 0 90 $X=58420 $Y=27110
X299 25 M2_M1_CDNS_9 $T=58670 31610 0 90 $X=58420 $Y=31530
X300 25 M2_M1_CDNS_9 $T=58670 38930 0 90 $X=58420 $Y=38850
X301 25 M2_M1_CDNS_9 $T=58670 46250 0 90 $X=58420 $Y=46170
X302 25 M2_M1_CDNS_9 $T=58670 53570 0 90 $X=58420 $Y=53490
X303 69 M2_M1_CDNS_9 $T=59660 13790 0 0 $X=59580 $Y=13540
X304 63 M2_M1_CDNS_9 $T=59660 21120 0 0 $X=59580 $Y=20870
X305 68 M2_M1_CDNS_9 $T=59660 28470 0 0 $X=59580 $Y=28220
X306 68 M5_M4_CDNS_10 $T=31030 6520 0 0 $X=30950 $Y=6390
X307 55 M5_M4_CDNS_10 $T=33450 34810 0 0 $X=33370 $Y=34680
X308 55 M5_M4_CDNS_10 $T=34490 38940 0 0 $X=34410 $Y=38810
X309 55 M5_M4_CDNS_10 $T=35140 50450 0 0 $X=35060 $Y=50320
X310 56 M5_M4_CDNS_10 $T=35270 23970 0 0 $X=35190 $Y=23840
X311 55 M5_M4_CDNS_10 $T=35630 42220 0 0 $X=35550 $Y=42090
X312 68 M5_M4_CDNS_10 $T=35740 16590 0 0 $X=35660 $Y=16460
X313 54 M5_M4_CDNS_10 $T=36550 34300 0 0 $X=36470 $Y=34170
X314 47 M5_M4_CDNS_10 $T=36920 33010 0 0 $X=36840 $Y=32880
X315 63 M5_M4_CDNS_10 $T=37650 13930 0 0 $X=37570 $Y=13800
X316 61 M5_M4_CDNS_10 $T=37800 9740 0 0 $X=37720 $Y=9610
X317 69 M5_M4_CDNS_10 $T=38000 8190 0 0 $X=37920 $Y=8060
X318 64 M5_M4_CDNS_10 $T=38690 18860 0 90 $X=38560 $Y=18780
X319 62 M5_M4_CDNS_10 $T=38750 26290 0 90 $X=38620 $Y=26210
X320 64 M5_M4_CDNS_10 $T=40200 18860 0 90 $X=40070 $Y=18780
X321 69 M5_M4_CDNS_10 $T=40300 8620 0 90 $X=40170 $Y=8540
X322 71 M5_M4_CDNS_10 $T=48360 8140 0 0 $X=48280 $Y=8010
X323 71 M5_M4_CDNS_10 $T=50330 8160 0 0 $X=50250 $Y=8030
X324 47 M5_M4_CDNS_10 $T=50340 37430 0 0 $X=50260 $Y=37300
X325 72 M3_M2_CDNS_11 $T=15150 34320 0 0 $X=15070 $Y=34070
X326 73 M3_M2_CDNS_11 $T=30360 48950 0 0 $X=30280 $Y=48700
X327 51 M3_M2_CDNS_11 $T=30540 30290 0 90 $X=30290 $Y=30210
X328 65 M3_M2_CDNS_11 $T=30920 28440 0 90 $X=30670 $Y=28360
X329 65 M3_M2_CDNS_11 $T=30920 23090 0 0 $X=30840 $Y=22840
X330 51 M3_M2_CDNS_11 $T=30960 32190 0 0 $X=30880 $Y=31940
X331 60 M3_M2_CDNS_11 $T=34240 15510 0 0 $X=34160 $Y=15260
X332 62 M3_M2_CDNS_11 $T=36070 26280 0 0 $X=35990 $Y=26030
X333 51 M3_M2_CDNS_11 $T=36600 41550 0 0 $X=36520 $Y=41300
X334 56 M3_M2_CDNS_11 $T=37800 29000 0 0 $X=37720 $Y=28750
X335 70 M3_M2_CDNS_11 $T=40600 12040 0 0 $X=40520 $Y=11790
X336 71 M3_M2_CDNS_11 $T=41660 8130 0 0 $X=41580 $Y=7880
X337 69 M3_M2_CDNS_11 $T=43120 8620 0 0 $X=43040 $Y=8370
X338 7 M3_M2_CDNS_11 $T=45720 13840 0 0 $X=45640 $Y=13590
X339 7 M3_M2_CDNS_11 $T=47400 30300 0 0 $X=47320 $Y=30050
X340 47 M3_M2_CDNS_11 $T=50830 40760 0 90 $X=50580 $Y=40680
X341 25 M3_M2_CDNS_11 $T=58260 1650 0 0 $X=58180 $Y=1400
X342 5 M4_M3_CDNS_12 $T=1340 55390 0 0 $X=1260 $Y=55140
X343 5 M4_M3_CDNS_12 $T=3450 61970 0 0 $X=3370 $Y=61720
X344 5 M4_M3_CDNS_12 $T=9870 69280 0 0 $X=9790 $Y=69030
X345 50 M4_M3_CDNS_12 $T=14700 34240 0 0 $X=14620 $Y=33990
X346 72 M4_M3_CDNS_12 $T=15150 34320 0 0 $X=15070 $Y=34070
X347 67 M4_M3_CDNS_12 $T=28040 20980 0 0 $X=27960 $Y=20730
X348 73 M4_M3_CDNS_12 $T=30360 48950 0 0 $X=30280 $Y=48700
X349 51 M4_M3_CDNS_12 $T=30540 30290 0 90 $X=30290 $Y=30210
X350 65 M4_M3_CDNS_12 $T=30920 28440 0 90 $X=30670 $Y=28360
X351 65 M4_M3_CDNS_12 $T=30920 23090 0 0 $X=30840 $Y=22840
X352 51 M4_M3_CDNS_12 $T=30960 32190 0 0 $X=30880 $Y=31940
X353 60 M4_M3_CDNS_12 $T=34240 15510 0 0 $X=34160 $Y=15260
X354 62 M4_M3_CDNS_12 $T=36070 26280 0 0 $X=35990 $Y=26030
X355 51 M4_M3_CDNS_12 $T=36600 41550 0 0 $X=36520 $Y=41300
X356 49 M4_M3_CDNS_12 $T=37620 30320 0 0 $X=37540 $Y=30070
X357 56 M4_M3_CDNS_12 $T=37800 29000 0 0 $X=37720 $Y=28750
X358 51 M4_M3_CDNS_12 $T=38820 45300 0 0 $X=38740 $Y=45050
X359 70 M4_M3_CDNS_12 $T=40600 12040 0 0 $X=40520 $Y=11790
X360 70 M4_M3_CDNS_12 $T=40600 13810 0 0 $X=40520 $Y=13560
X361 71 M4_M3_CDNS_12 $T=41660 8130 0 0 $X=41580 $Y=7880
X362 69 M4_M3_CDNS_12 $T=43120 8620 0 0 $X=43040 $Y=8370
X363 7 M4_M3_CDNS_12 $T=45720 13840 0 0 $X=45640 $Y=13590
X364 7 M4_M3_CDNS_12 $T=46890 13630 0 0 $X=46810 $Y=13380
X365 7 M4_M3_CDNS_12 $T=46900 20740 0 0 $X=46820 $Y=20490
X366 7 M4_M3_CDNS_12 $T=46910 28080 0 0 $X=46830 $Y=27830
X367 5 M4_M3_CDNS_12 $T=49180 4060 0 0 $X=49100 $Y=3810
X368 5 M4_M3_CDNS_12 $T=49180 11470 0 0 $X=49100 $Y=11220
X369 5 M4_M3_CDNS_12 $T=49180 18800 0 0 $X=49100 $Y=18550
X370 5 M4_M3_CDNS_12 $T=49180 26120 0 0 $X=49100 $Y=25870
X371 5 M4_M3_CDNS_12 $T=49180 33430 0 0 $X=49100 $Y=33180
X372 5 M4_M3_CDNS_12 $T=49180 40820 0 0 $X=49100 $Y=40570
X373 5 M4_M3_CDNS_12 $T=49180 48070 0 0 $X=49100 $Y=47820
X374 5 M4_M3_CDNS_12 $T=49180 54710 0 0 $X=49100 $Y=54460
X375 47 M4_M3_CDNS_12 $T=50830 40760 0 90 $X=50580 $Y=40680
X376 25 M4_M3_CDNS_12 $T=58260 1650 0 0 $X=58180 $Y=1400
X377 25 M4_M3_CDNS_12 $T=58670 9650 0 90 $X=58420 $Y=9570
X378 25 M4_M3_CDNS_12 $T=58670 12550 0 90 $X=58420 $Y=12470
X379 25 M4_M3_CDNS_12 $T=58670 16970 0 90 $X=58420 $Y=16890
X380 25 M4_M3_CDNS_12 $T=58670 19870 0 90 $X=58420 $Y=19790
X381 25 M4_M3_CDNS_12 $T=58670 24290 0 90 $X=58420 $Y=24210
X382 25 M4_M3_CDNS_12 $T=58670 27190 0 90 $X=58420 $Y=27110
X383 25 M4_M3_CDNS_12 $T=58670 31610 0 90 $X=58420 $Y=31530
X384 25 M4_M3_CDNS_12 $T=58670 38930 0 90 $X=58420 $Y=38850
X385 25 M4_M3_CDNS_12 $T=58670 46250 0 90 $X=58420 $Y=46170
X386 25 M4_M3_CDNS_12 $T=58670 53570 0 90 $X=58420 $Y=53490
X387 50 M4_M3_CDNS_13 $T=13710 9140 0 0 $X=13630 $Y=9010
X388 50 M4_M3_CDNS_13 $T=13710 17480 0 0 $X=13630 $Y=17350
X389 50 M4_M3_CDNS_13 $T=13710 19960 0 0 $X=13630 $Y=19830
X390 72 M4_M3_CDNS_13 $T=14090 21060 0 0 $X=14010 $Y=20930
X391 48 M4_M3_CDNS_13 $T=24590 43490 0 0 $X=24510 $Y=43360
X392 73 M4_M3_CDNS_13 $T=28000 27530 0 0 $X=27920 $Y=27400
X393 48 M4_M3_CDNS_13 $T=28120 30940 0 0 $X=28040 $Y=30810
X394 63 M4_M3_CDNS_13 $T=30320 6550 0 0 $X=30240 $Y=6420
X395 68 M4_M3_CDNS_13 $T=31030 8560 0 90 $X=30900 $Y=8480
X396 61 M4_M3_CDNS_13 $T=34270 8400 0 0 $X=34190 $Y=8270
X397 49 M4_M3_CDNS_13 $T=34570 23190 0 0 $X=34490 $Y=23060
X398 68 M4_M3_CDNS_13 $T=34690 12200 0 0 $X=34610 $Y=12070
X399 47 M4_M3_CDNS_13 $T=36100 30140 0 0 $X=36020 $Y=30010
X400 54 M4_M3_CDNS_13 $T=36540 37650 0 90 $X=36410 $Y=37570
X401 60 M4_M3_CDNS_13 $T=37250 15560 0 0 $X=37170 $Y=15430
X402 67 M4_M3_CDNS_13 $T=37310 22870 0 0 $X=37230 $Y=22740
X403 66 M4_M3_CDNS_13 $T=37550 19040 0 0 $X=37470 $Y=18910
X404 66 M4_M3_CDNS_13 $T=37670 21700 0 0 $X=37590 $Y=21570
X405 64 M4_M3_CDNS_13 $T=38370 9550 0 0 $X=38290 $Y=9420
X406 64 M4_M3_CDNS_13 $T=40710 21060 0 0 $X=40630 $Y=20930
X407 69 M4_M3_CDNS_13 $T=41120 2720 0 0 $X=41040 $Y=2590
X408 7 M4_M3_CDNS_13 $T=47400 30300 0 0 $X=47320 $Y=30170
X409 6 M4_M3_CDNS_13 $T=48170 14160 0 0 $X=48090 $Y=14030
X410 6 M4_M3_CDNS_13 $T=48170 17210 0 0 $X=48090 $Y=17080
X411 71 M4_M3_CDNS_13 $T=50910 13780 0 0 $X=50830 $Y=13650
X412 6 M1_PO_CDNS_14 $T=1860 60810 0 0 $X=1760 $Y=60560
X413 6 M1_PO_CDNS_14 $T=1870 68120 0 0 $X=1770 $Y=67870
X414 4 M1_PO_CDNS_14 $T=2350 44590 0 90 $X=2100 $Y=44490
X415 3 M1_PO_CDNS_14 $T=3900 48300 0 90 $X=3650 $Y=48200
X416 2 M1_PO_CDNS_14 $T=3940 58210 0 90 $X=3690 $Y=58110
X417 11 M1_PO_CDNS_14 $T=6840 58120 0 90 $X=6590 $Y=58020
X418 6 M1_PO_CDNS_14 $T=12100 60800 0 0 $X=12000 $Y=60550
X419 6 M1_PO_CDNS_14 $T=12100 68120 0 0 $X=12000 $Y=67870
X420 6 M1_PO_CDNS_14 $T=22340 68120 0 0 $X=22240 $Y=67870
X421 6 M1_PO_CDNS_14 $T=22350 60800 0 0 $X=22250 $Y=60550
X422 6 M1_PO_CDNS_14 $T=32580 60800 0 0 $X=32480 $Y=60550
X423 6 M1_PO_CDNS_14 $T=32580 68120 0 0 $X=32480 $Y=67870
X424 68 M1_PO_CDNS_14 $T=33670 6150 0 90 $X=33420 $Y=6050
X425 6 M1_PO_CDNS_14 $T=40360 10220 0 90 $X=40110 $Y=10120
X426 6 M1_PO_CDNS_14 $T=40340 24940 0 0 $X=40240 $Y=24690
X427 6 M1_PO_CDNS_14 $T=40370 17590 0 0 $X=40270 $Y=17340
X428 7 M1_PO_CDNS_14 $T=46890 13630 0 0 $X=46790 $Y=13380
X429 7 M1_PO_CDNS_14 $T=46900 20740 0 0 $X=46800 $Y=20490
X430 7 M1_PO_CDNS_14 $T=46910 28080 0 0 $X=46810 $Y=27830
X431 6 M1_PO_CDNS_14 $T=47620 54480 0 90 $X=47370 $Y=54380
X432 6 M1_PO_CDNS_14 $T=47800 38230 0 90 $X=47550 $Y=38130
X433 6 M1_PO_CDNS_14 $T=47870 10240 0 0 $X=47770 $Y=9990
X434 6 M1_PO_CDNS_14 $T=47980 9490 0 0 $X=47880 $Y=9240
X435 6 M1_PO_CDNS_14 $T=48260 51950 0 90 $X=48010 $Y=51850
X436 6 M1_PO_CDNS_14 $T=48260 45130 0 0 $X=48160 $Y=44880
X437 6 M1_PO_CDNS_14 $T=48690 16910 0 0 $X=48590 $Y=16660
X438 6 M1_PO_CDNS_14 $T=48860 24230 0 0 $X=48760 $Y=23980
X439 6 M1_PO_CDNS_14 $T=48880 2280 0 0 $X=48780 $Y=2030
X440 6 M1_PO_CDNS_15 $T=47780 31470 0 0 $X=47680 $Y=31220
X441 7 M1_PO_CDNS_16 $T=47950 48930 0 0 $X=47850 $Y=48810
X442 6 M2_M1_CDNS_17 $T=47780 31470 0 0 $X=47700 $Y=31220
X443 1 5 2 3 4 10 15 14 11 50
+ 16 46 72 48 53 65 51 73 251 260
+ 231 228 214 224 218 288 249 250 253 313
+ 314 307 275 219 266 278 216 289 290 277
+ 293 318 232 279 296 317 300 262 316 261 multiplier $T=1090 33260 0 0 $X=750 $Y=33040
X444 63 8 10 5 9 65 48 68 61 58
+ 56 49 54 55 73 51 72 57 53 50
+ 46 64 69 19 59 67 47 52 66 71
+ 60 62 70 74 95 112 111 110 109 115
+ 114 121 120 119 118 103 102 105 104 141
+ 211 107 106 97 96 99 98 101 100 108
+ 113 130 139 140 158 159 176 185 190 191
+ 194 212 213 760 761 762 763 10badder $T=-50390 53780 1 0 $X=-110 $Y=0
X445 10 7 5 6 1 12 90 86 91 87
+ 506 88 508 84 85 89 92 ph1p3_MSDFF $T=1140 62320 0 0 $X=1140 $Y=58560
X446 10 7 5 6 2 13 81 77 82 78
+ 503 79 505 75 76 80 83 ph1p3_MSDFF $T=1140 69640 0 0 $X=1140 $Y=65880
X447 10 7 5 6 15 18 345 341 346 342
+ 692 343 694 339 340 344 347 ph1p3_MSDFF $T=11380 62320 0 0 $X=11380 $Y=58560
X448 10 7 5 6 11 17 336 332 337 333
+ 689 334 691 330 331 335 338 ph1p3_MSDFF $T=11380 69640 0 0 $X=11380 $Y=65880
X449 10 7 5 6 14 21 363 359 364 360
+ 698 361 700 357 358 362 365 ph1p3_MSDFF $T=21620 62320 0 0 $X=21620 $Y=58560
X450 10 7 5 6 3 20 354 350 355 351
+ 695 352 697 348 349 353 356 ph1p3_MSDFF $T=21620 69640 0 0 $X=21620 $Y=65880
X451 10 7 5 6 16 22 381 377 382 378
+ 704 379 706 375 376 380 383 ph1p3_MSDFF $T=31860 62320 0 0 $X=31860 $Y=58560
X452 10 7 5 6 4 23 372 368 373 369
+ 701 370 703 366 367 371 374 ph1p3_MSDFF $T=31860 69640 0 0 $X=31860 $Y=65880
X453 10 7 5 6 70 69 408 404 409 405
+ 713 406 715 402 403 407 410 ph1p3_MSDFF $T=37920 11080 0 0 $X=37920 $Y=7320
X454 10 7 5 6 64 63 399 395 400 396
+ 710 397 712 393 394 398 401 ph1p3_MSDFF $T=37920 18400 0 0 $X=37920 $Y=14640
X455 10 7 5 6 66 68 390 386 391 387
+ 707 388 709 384 385 389 392 ph1p3_MSDFF $T=37920 25720 0 0 $X=37920 $Y=21960
X456 10 7 5 6 24 25 480 476 481 477
+ 737 478 739 474 475 479 482 ph1p3_MSDFF $T=48160 3760 0 0 $X=48160 $Y=0
X457 10 7 5 6 71 61 471 467 472 468
+ 734 469 736 465 466 470 473 ph1p3_MSDFF $T=48160 11080 0 0 $X=48160 $Y=7320
X458 10 7 5 6 60 58 462 458 463 459
+ 731 460 733 456 457 461 464 ph1p3_MSDFF $T=48160 18400 0 0 $X=48160 $Y=14640
X459 10 7 5 6 62 57 453 449 454 450
+ 728 451 730 447 448 452 455 ph1p3_MSDFF $T=48160 25720 0 0 $X=48160 $Y=21960
X460 10 7 5 6 67 56 444 440 445 441
+ 725 442 727 438 439 443 446 ph1p3_MSDFF $T=48160 33040 0 0 $X=48160 $Y=29280
X461 10 7 5 6 47 49 435 431 436 432
+ 722 433 724 429 430 434 437 ph1p3_MSDFF $T=48160 40360 0 0 $X=48160 $Y=36600
X462 10 7 5 6 52 54 426 422 427 423
+ 719 424 721 420 421 425 428 ph1p3_MSDFF $T=48160 47680 0 0 $X=48160 $Y=43920
X463 10 7 5 6 59 55 417 413 418 414
+ 716 415 718 411 412 416 419 ph1p3_MSDFF $T=48160 55000 0 0 $X=48160 $Y=51240
X464 10 5 cellTmpl_CDNS_49 $T=47620 54900 1 0 $X=47500 $Y=51240
X465 25 61 10 5 36 34 501 502 758 759
+ 788 789 MUX_2to1___2X_ph2p2 $T=58160 11120 1 0 $X=58160 $Y=7320
X466 25 69 10 5 37 29 499 500 756 757
+ 786 787 MUX_2to1___2X_ph2p2 $T=58160 11080 0 0 $X=58160 $Y=11080
X467 25 58 10 5 38 26 497 498 754 755
+ 784 785 MUX_2to1___2X_ph2p2 $T=58160 18440 1 0 $X=58160 $Y=14640
X468 25 63 10 5 39 31 495 496 752 753
+ 782 783 MUX_2to1___2X_ph2p2 $T=58160 18400 0 0 $X=58160 $Y=18400
X469 25 57 10 5 40 32 493 494 750 751
+ 780 781 MUX_2to1___2X_ph2p2 $T=58160 25760 1 0 $X=58160 $Y=21960
X470 25 68 10 5 41 35 491 492 748 749
+ 778 779 MUX_2to1___2X_ph2p2 $T=58160 25720 0 0 $X=58160 $Y=25720
X471 25 56 10 5 42 28 489 490 746 747
+ 776 777 MUX_2to1___2X_ph2p2 $T=58160 33080 1 0 $X=58160 $Y=29280
X472 25 49 10 5 43 33 487 488 744 745
+ 774 775 MUX_2to1___2X_ph2p2 $T=58160 40400 1 0 $X=58160 $Y=36600
X473 25 54 10 5 44 30 485 486 742 743
+ 772 773 MUX_2to1___2X_ph2p2 $T=58160 47720 1 0 $X=58160 $Y=43920
X474 25 55 10 5 45 27 483 484 740 741
+ 770 771 MUX_2to1___2X_ph2p2 $T=58160 55040 1 0 $X=58160 $Y=51240
M0 87 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=59450 $dt=1
M1 90 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=64750 $dt=1
M2 78 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=1920 $Y=66770 $dt=1
M3 84 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3250 $Y=64780 $dt=1
M4 85 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=59420 $dt=1
M5 76 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=4250 $Y=66740 $dt=1
M6 86 7 1 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4430 $Y=64780 $dt=1
M7 91 7 506 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=59660 $dt=1
M8 82 7 503 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=5430 $Y=66980 $dt=1
M9 88 86 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=5630 $Y=64690 $dt=1
M10 506 12 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=59450 $dt=1
M11 503 13 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=6720 $Y=66770 $dt=1
M12 88 87 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=6870 $Y=64700 $dt=1
M13 89 90 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=59420 $dt=1
M14 80 81 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=8050 $Y=66740 $dt=1
M15 508 88 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8120 $Y=64750 $dt=1
M16 91 90 88 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=59660 $dt=1
M17 82 81 79 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=9230 $Y=66980 $dt=1
M18 92 90 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9450 $Y=64780 $dt=1
M19 12 91 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=59450 $dt=1
M20 13 82 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=10520 $Y=66770 $dt=1
M21 86 90 508 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=10630 $Y=64780 $dt=1
M22 342 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=59450 $dt=1
M23 345 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=64750 $dt=1
M24 333 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12160 $Y=66770 $dt=1
M25 339 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13490 $Y=64780 $dt=1
M26 340 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=59420 $dt=1
M27 331 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=14490 $Y=66740 $dt=1
M28 341 7 15 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=14670 $Y=64780 $dt=1
M29 346 7 692 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=59660 $dt=1
M30 337 7 689 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15670 $Y=66980 $dt=1
M31 343 341 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=15870 $Y=64690 $dt=1
M32 692 18 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=59450 $dt=1
M33 689 17 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=16960 $Y=66770 $dt=1
M34 343 342 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17110 $Y=64700 $dt=1
M35 344 345 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=59420 $dt=1
M36 335 336 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=18290 $Y=66740 $dt=1
M37 694 343 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18360 $Y=64750 $dt=1
M38 346 345 343 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=59660 $dt=1
M39 337 336 334 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=19470 $Y=66980 $dt=1
M40 347 345 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=19690 $Y=64780 $dt=1
M41 18 346 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=59450 $dt=1
M42 17 337 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=20760 $Y=66770 $dt=1
M43 341 345 694 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=20870 $Y=64780 $dt=1
M44 360 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=59450 $dt=1
M45 363 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=64750 $dt=1
M46 351 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22400 $Y=66770 $dt=1
M47 357 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=23730 $Y=64780 $dt=1
M48 358 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=59420 $dt=1
M49 349 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24730 $Y=66740 $dt=1
M50 359 7 14 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=24910 $Y=64780 $dt=1
M51 364 7 698 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=59660 $dt=1
M52 355 7 695 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25910 $Y=66980 $dt=1
M53 361 359 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26110 $Y=64690 $dt=1
M54 698 21 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=59450 $dt=1
M55 695 20 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=27200 $Y=66770 $dt=1
M56 361 360 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27350 $Y=64700 $dt=1
M57 362 363 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=59420 $dt=1
M58 353 354 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=28530 $Y=66740 $dt=1
M59 700 361 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28600 $Y=64750 $dt=1
M60 364 363 361 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=59660 $dt=1
M61 355 354 352 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=29710 $Y=66980 $dt=1
M62 365 363 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=29930 $Y=64780 $dt=1
M63 21 364 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=59450 $dt=1
M64 20 355 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=31000 $Y=66770 $dt=1
M65 359 363 700 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31110 $Y=64780 $dt=1
M66 378 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=59450 $dt=1
M67 381 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=64750 $dt=1
M68 369 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=32640 $Y=66770 $dt=1
M69 375 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=33970 $Y=64780 $dt=1
M70 376 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=59420 $dt=1
M71 367 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34970 $Y=66740 $dt=1
M72 377 7 16 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35150 $Y=64780 $dt=1
M73 382 7 704 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=59660 $dt=1
M74 373 7 701 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=36150 $Y=66980 $dt=1
M75 379 377 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36350 $Y=64690 $dt=1
M76 704 22 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=37440 $Y=59450 $dt=1
M77 701 23 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=37440 $Y=66770 $dt=1
M78 379 378 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37590 $Y=64700 $dt=1
M79 405 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=8210 $dt=1
M80 408 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=13510 $dt=1
M81 396 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=15530 $dt=1
M82 399 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=20830 $dt=1
M83 387 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=38700 $Y=22850 $dt=1
M84 390 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=38700 $Y=28150 $dt=1
M85 380 381 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=38770 $Y=59420 $dt=1
M86 371 372 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=38770 $Y=66740 $dt=1
M87 706 379 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=38840 $Y=64750 $dt=1
M88 382 381 379 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=39950 $Y=59660 $dt=1
M89 373 372 370 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=39950 $Y=66980 $dt=1
M90 402 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=13540 $dt=1
M91 393 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=40030 $Y=20860 $dt=1
M92 384 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=40030 $Y=28180 $dt=1
M93 383 381 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40170 $Y=64780 $dt=1
M94 403 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=41030 $Y=8180 $dt=1
M95 394 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=15500 $dt=1
M96 385 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=41030 $Y=22820 $dt=1
M97 404 7 70 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=13540 $dt=1
M98 395 7 64 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=41210 $Y=20860 $dt=1
M99 386 7 66 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=41210 $Y=28180 $dt=1
M100 22 382 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=41240 $Y=59450 $dt=1
M101 23 373 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.2497 scb=0.0129015 scc=0.000236549 $X=41240 $Y=66770 $dt=1
M102 377 381 706 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41350 $Y=64780 $dt=1
M103 409 7 713 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=42210 $Y=8420 $dt=1
M104 400 7 710 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=15740 $dt=1
M105 391 7 707 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=42210 $Y=23060 $dt=1
M106 406 404 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=13450 $dt=1
M107 397 395 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=42410 $Y=20770 $dt=1
M108 388 386 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=42410 $Y=28090 $dt=1
M109 713 69 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=43500 $Y=8210 $dt=1
M110 710 63 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=15530 $dt=1
M111 707 68 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=43500 $Y=22850 $dt=1
M112 406 405 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=13460 $dt=1
M113 397 396 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=43650 $Y=20780 $dt=1
M114 388 387 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=43650 $Y=28100 $dt=1
M115 407 408 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=44830 $Y=8180 $dt=1
M116 398 399 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=15500 $dt=1
M117 389 390 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=44830 $Y=22820 $dt=1
M118 715 406 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=13510 $dt=1
M119 712 397 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=44900 $Y=20830 $dt=1
M120 709 388 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=44900 $Y=28150 $dt=1
M121 409 408 406 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=46010 $Y=8420 $dt=1
M122 400 399 397 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=15740 $dt=1
M123 391 390 388 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=46010 $Y=23060 $dt=1
M124 410 408 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=13540 $dt=1
M125 401 399 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=46230 $Y=20860 $dt=1
M126 392 390 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=46230 $Y=28180 $dt=1
M127 69 409 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=47300 $Y=8210 $dt=1
M128 63 400 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=15530 $dt=1
M129 68 391 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=47300 $Y=22850 $dt=1
M130 404 408 715 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=13540 $dt=1
M131 395 399 712 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=47410 $Y=20860 $dt=1
M132 386 390 709 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=47410 $Y=28180 $dt=1
M133 477 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=890 $dt=1
M134 480 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=6190 $dt=1
M135 468 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=8210 $dt=1
M136 471 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=13510 $dt=1
M137 459 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=15530 $dt=1
M138 462 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=20830 $dt=1
M139 450 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=22850 $dt=1
M140 453 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=28150 $dt=1
M141 441 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=30170 $dt=1
M142 444 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=35470 $dt=1
M143 432 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=37490 $dt=1
M144 435 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=42790 $dt=1
M145 423 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=44810 $dt=1
M146 426 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=48940 $Y=50110 $dt=1
M147 414 6 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=48940 $Y=52130 $dt=1
M148 417 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=48940 $Y=57430 $dt=1
M149 474 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=6220 $dt=1
M150 465 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=13540 $dt=1
M151 456 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=20860 $dt=1
M152 447 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=28180 $dt=1
M153 438 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=35500 $dt=1
M154 429 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=42820 $dt=1
M155 420 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=50270 $Y=50140 $dt=1
M156 411 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=50270 $Y=57460 $dt=1
M157 475 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=51270 $Y=860 $dt=1
M158 466 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=8180 $dt=1
M159 457 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=15500 $dt=1
M160 448 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=22820 $dt=1
M161 439 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=30140 $dt=1
M162 430 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=37460 $dt=1
M163 421 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=44780 $dt=1
M164 412 7 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=51270 $Y=52100 $dt=1
M165 476 7 24 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=6220 $dt=1
M166 467 7 71 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=13540 $dt=1
M167 458 7 60 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=20860 $dt=1
M168 449 7 62 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=28180 $dt=1
M169 440 7 67 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=35500 $dt=1
M170 431 7 47 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=42820 $dt=1
M171 422 7 52 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=51450 $Y=50140 $dt=1
M172 413 7 59 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=51450 $Y=57460 $dt=1
M173 481 7 737 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=52450 $Y=1100 $dt=1
M174 472 7 734 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=8420 $dt=1
M175 463 7 731 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=15740 $dt=1
M176 454 7 728 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=23060 $dt=1
M177 445 7 725 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=30380 $dt=1
M178 436 7 722 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=37700 $dt=1
M179 427 7 719 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=45020 $dt=1
M180 418 7 716 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=52450 $Y=52340 $dt=1
M181 478 476 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=6130 $dt=1
M182 469 467 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=13450 $dt=1
M183 460 458 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=20770 $dt=1
M184 451 449 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=28090 $dt=1
M185 442 440 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=35410 $dt=1
M186 433 431 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=42730 $dt=1
M187 424 422 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=52650 $Y=50050 $dt=1
M188 415 413 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=52650 $Y=57370 $dt=1
M189 737 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=53740 $Y=890 $dt=1
M190 734 61 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=8210 $dt=1
M191 731 58 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=15530 $dt=1
M192 728 57 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=22850 $dt=1
M193 725 56 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=30170 $dt=1
M194 722 49 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=37490 $dt=1
M195 719 54 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=44810 $dt=1
M196 716 55 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=53740 $Y=52130 $dt=1
M197 478 477 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=6140 $dt=1
M198 469 468 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=13460 $dt=1
M199 460 459 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=20780 $dt=1
M200 451 450 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=28100 $dt=1
M201 442 441 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=35420 $dt=1
M202 433 432 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=42740 $dt=1
M203 424 423 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=53890 $Y=50060 $dt=1
M204 415 414 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=53890 $Y=57380 $dt=1
M205 479 480 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=55070 $Y=860 $dt=1
M206 470 471 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=8180 $dt=1
M207 461 462 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=15500 $dt=1
M208 452 453 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=22820 $dt=1
M209 443 444 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=30140 $dt=1
M210 434 435 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=37460 $dt=1
M211 425 426 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=44780 $dt=1
M212 416 417 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=55070 $Y=52100 $dt=1
M213 739 478 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=6190 $dt=1
M214 736 469 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=13510 $dt=1
M215 733 460 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=20830 $dt=1
M216 730 451 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=28150 $dt=1
M217 727 442 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=35470 $dt=1
M218 724 433 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=42790 $dt=1
M219 721 424 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=55140 $Y=50110 $dt=1
M220 718 415 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=55140 $Y=57430 $dt=1
M221 481 480 478 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=56250 $Y=1100 $dt=1
M222 472 471 469 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=8420 $dt=1
M223 463 462 460 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=15740 $dt=1
M224 454 453 451 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=23060 $dt=1
M225 445 444 442 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=30380 $dt=1
M226 436 435 433 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=37700 $dt=1
M227 427 426 424 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=45020 $dt=1
M228 418 417 415 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=56250 $Y=52340 $dt=1
M229 482 480 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=6220 $dt=1
M230 473 471 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=13540 $dt=1
M231 464 462 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=20860 $dt=1
M232 455 453 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=56470 $Y=28180 $dt=1
M233 446 444 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=35500 $dt=1
M234 437 435 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=42820 $dt=1
M235 428 426 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=56470 $Y=50140 $dt=1
M236 419 417 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=56470 $Y=57460 $dt=1
M237 25 481 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.7239 scb=0.0151885 scc=0.000250442 $X=57540 $Y=890 $dt=1
M238 61 472 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=8210 $dt=1
M239 58 463 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=15530 $dt=1
M240 57 454 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=22850 $dt=1
M241 56 445 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=30170 $dt=1
M242 49 436 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=37490 $dt=1
M243 54 427 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=44810 $dt=1
M244 55 418 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=57540 $Y=52130 $dt=1
M245 476 480 739 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=6220 $dt=1
M246 467 471 736 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=13540 $dt=1
M247 458 462 733 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=20860 $dt=1
M248 449 453 730 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=57650 $Y=28180 $dt=1
M249 440 444 727 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=35500 $dt=1
M250 431 435 724 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=42820 $dt=1
M251 422 426 721 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=57650 $Y=50140 $dt=1
M252 413 417 718 10 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=57650 $Y=57460 $dt=1
M253 501 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=8270 $dt=1
M254 499 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=13450 $dt=1
M255 497 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=15590 $dt=1
M256 495 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=20770 $dt=1
M257 493 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=22910 $dt=1
M258 491 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=28090 $dt=1
M259 489 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=59090 $Y=30230 $dt=1
M260 487 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=37550 $dt=1
M261 485 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=44870 $dt=1
M262 483 25 10 10 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=59090 $Y=52190 $dt=1
M263 788 61 502 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=8060 $dt=1
M264 786 69 500 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=13180 $dt=1
M265 784 58 498 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=15380 $dt=1
M266 782 63 496 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=20500 $dt=1
M267 780 57 494 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=22700 $dt=1
M268 778 68 492 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=27820 $dt=1
M269 776 56 490 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60120 $Y=30020 $dt=1
M270 774 49 488 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=37340 $dt=1
M271 772 54 486 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=44660 $dt=1
M272 770 55 484 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60120 $Y=51980 $dt=1
M273 10 25 788 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=8060 $dt=1
M274 10 25 786 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=13180 $dt=1
M275 10 25 784 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=15380 $dt=1
M276 10 25 782 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=20500 $dt=1
M277 10 25 780 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=22700 $dt=1
M278 10 25 778 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=27820 $dt=1
M279 10 25 776 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=60330 $Y=30020 $dt=1
M280 10 25 774 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=37340 $dt=1
M281 10 25 772 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=44660 $dt=1
M282 10 25 770 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=60330 $Y=51980 $dt=1
M283 789 501 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=8130 $dt=1
M284 787 499 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=13110 $dt=1
M285 785 497 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=15450 $dt=1
M286 783 495 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=20430 $dt=1
M287 781 493 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=22770 $dt=1
M288 779 491 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=27750 $dt=1
M289 777 489 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61500 $Y=30090 $dt=1
M290 775 487 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=37410 $dt=1
M291 773 485 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=44730 $dt=1
M292 771 483 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=2.88e-14 AS=6.72e-14 PD=1.08e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=2.45e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61500 $Y=52050 $dt=1
M293 502 36 789 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=8130 $dt=1
M294 500 37 787 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=13110 $dt=1
M295 498 38 785 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=15450 $dt=1
M296 496 39 783 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=20430 $dt=1
M297 494 40 781 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=22770 $dt=1
M298 492 41 779 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=27750 $dt=1
M299 490 42 777 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=15.8127 scb=0.0131685 scc=0.00149596 $X=61710 $Y=30090 $dt=1
M300 488 43 775 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=37410 $dt=1
M301 486 44 773 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=44730 $dt=1
M302 484 45 771 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=2.88e-14 PD=1.24e-06 PS=1.08e-06 fw=4.8e-07 sa=2.45e-07 sb=1.4e-07 sca=17.927 scb=0.0149618 scc=0.00151035 $X=61710 $Y=52050 $dt=1
M303 34 502 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=8120 $dt=1
M304 29 500 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=13120 $dt=1
M305 26 498 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=15440 $dt=1
M306 31 496 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=20440 $dt=1
M307 32 494 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=22760 $dt=1
M308 35 492 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=27760 $dt=1
M309 28 490 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=19.9967 scb=0.019222 scc=0.00149353 $X=62920 $Y=30080 $dt=1
M310 33 488 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=37400 $dt=1
M311 30 486 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=44720 $dt=1
M312 27 484 10 10 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=22.1619 scb=0.0210888 scc=0.00150925 $X=62920 $Y=52040 $dt=1
.ends ph2p2_processing_element

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph2p3_Matrix_vector_Multiplication              *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph2p3_Matrix_vector_Multiplication 1 2 3 4 5 6 7 8 9 10
+ 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30
+ 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50
+ 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70
+ 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90
+ 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126
** N=2678 EP=126 FDC=6648
X0 11 M3_M2_CDNS_1 $T=47980 58060 0 90 $X=47730 $Y=57980
X1 11 M3_M2_CDNS_1 $T=47980 131280 0 90 $X=47730 $Y=131200
X2 11 M3_M2_CDNS_1 $T=47980 204490 0 90 $X=47730 $Y=204410
X3 85 M3_M2_CDNS_1 $T=63820 31300 0 0 $X=63740 $Y=31050
X4 85 M3_M2_CDNS_1 $T=63820 71930 0 0 $X=63740 $Y=71680
X5 86 M3_M2_CDNS_1 $T=63820 104520 0 0 $X=63740 $Y=104270
X6 86 M3_M2_CDNS_1 $T=63820 145150 0 0 $X=63740 $Y=144900
X7 87 M3_M2_CDNS_1 $T=63820 177730 0 0 $X=63740 $Y=177480
X8 87 M3_M2_CDNS_1 $T=63820 218360 0 0 $X=63740 $Y=218110
X9 88 M3_M2_CDNS_1 $T=63850 23980 0 0 $X=63770 $Y=23730
X10 89 M3_M2_CDNS_1 $T=63850 97200 0 0 $X=63770 $Y=96950
X11 90 M3_M2_CDNS_1 $T=63850 170410 0 0 $X=63770 $Y=170160
X12 91 M3_M2_CDNS_1 $T=63890 27300 0 0 $X=63810 $Y=27050
X13 92 M3_M2_CDNS_1 $T=63890 100520 0 0 $X=63810 $Y=100270
X14 93 M3_M2_CDNS_1 $T=63890 173730 0 0 $X=63810 $Y=173480
X15 11 M2_M1_CDNS_2 $T=47980 58060 0 90 $X=47730 $Y=57980
X16 11 M2_M1_CDNS_2 $T=47980 131280 0 90 $X=47730 $Y=131200
X17 11 M2_M1_CDNS_2 $T=47980 204490 0 90 $X=47730 $Y=204410
X18 85 M2_M1_CDNS_2 $T=63820 31300 0 0 $X=63740 $Y=31050
X19 85 M2_M1_CDNS_2 $T=63820 71930 0 0 $X=63740 $Y=71680
X20 86 M2_M1_CDNS_2 $T=63820 104520 0 0 $X=63740 $Y=104270
X21 86 M2_M1_CDNS_2 $T=63820 145150 0 0 $X=63740 $Y=144900
X22 87 M2_M1_CDNS_2 $T=63820 177730 0 0 $X=63740 $Y=177480
X23 87 M2_M1_CDNS_2 $T=63820 218360 0 0 $X=63740 $Y=218110
X24 88 M2_M1_CDNS_2 $T=63850 23980 0 0 $X=63770 $Y=23730
X25 89 M2_M1_CDNS_2 $T=63850 97200 0 0 $X=63770 $Y=96950
X26 90 M2_M1_CDNS_2 $T=63850 170410 0 0 $X=63770 $Y=170160
X27 91 M2_M1_CDNS_2 $T=63890 27300 0 0 $X=63810 $Y=27050
X28 92 M2_M1_CDNS_2 $T=63890 100520 0 0 $X=63810 $Y=100270
X29 93 M2_M1_CDNS_2 $T=63890 173730 0 0 $X=63810 $Y=173480
X30 85 M4_M3_CDNS_3 $T=49120 82570 0 0 $X=49040 $Y=82320
X31 86 M4_M3_CDNS_3 $T=49120 155790 0 0 $X=49040 $Y=155540
X32 87 M4_M3_CDNS_3 $T=49120 229000 0 0 $X=49040 $Y=228750
X33 94 M4_M3_CDNS_3 $T=53160 72250 0 0 $X=53080 $Y=72000
X34 95 M4_M3_CDNS_3 $T=53160 145470 0 0 $X=53080 $Y=145220
X35 96 M4_M3_CDNS_3 $T=53160 218680 0 0 $X=53080 $Y=218430
X36 94 M4_M3_CDNS_3 $T=55950 72850 0 90 $X=55700 $Y=72770
X37 95 M4_M3_CDNS_3 $T=55950 146070 0 90 $X=55700 $Y=145990
X38 96 M4_M3_CDNS_3 $T=55950 219280 0 90 $X=55700 $Y=219200
X39 85 M5_M4_CDNS_5 $T=49120 82570 0 0 $X=49040 $Y=82320
X40 86 M5_M4_CDNS_5 $T=49120 155790 0 0 $X=49040 $Y=155540
X41 87 M5_M4_CDNS_5 $T=49120 229000 0 0 $X=49040 $Y=228750
X42 94 M5_M4_CDNS_5 $T=53160 72250 0 0 $X=53080 $Y=72000
X43 95 M5_M4_CDNS_5 $T=53160 145470 0 0 $X=53080 $Y=145220
X44 96 M5_M4_CDNS_5 $T=53160 218680 0 0 $X=53080 $Y=218430
X45 94 M5_M4_CDNS_5 $T=55950 72850 0 90 $X=55700 $Y=72770
X46 95 M5_M4_CDNS_5 $T=55950 146070 0 90 $X=55700 $Y=145990
X47 96 M5_M4_CDNS_5 $T=55950 219280 0 90 $X=55700 $Y=219200
X48 85 M5_M4_CDNS_5 $T=62740 103290 0 0 $X=62660 $Y=103040
X49 86 M5_M4_CDNS_5 $T=62740 176510 0 0 $X=62660 $Y=176260
X50 87 M5_M4_CDNS_5 $T=62740 249720 0 0 $X=62660 $Y=249470
X51 97 M5_M4_CDNS_5 $T=62750 87190 0 0 $X=62670 $Y=86940
X52 98 M5_M4_CDNS_5 $T=62750 160410 0 0 $X=62670 $Y=160160
X53 99 M5_M4_CDNS_5 $T=62750 233620 0 0 $X=62670 $Y=233370
X54 100 M5_M4_CDNS_5 $T=62760 88540 0 0 $X=62680 $Y=88290
X55 101 M5_M4_CDNS_5 $T=62760 94470 0 0 $X=62680 $Y=94220
X56 88 M5_M4_CDNS_5 $T=62760 95900 0 0 $X=62680 $Y=95650
X57 91 M5_M4_CDNS_5 $T=62760 101860 0 0 $X=62680 $Y=101610
X58 102 M5_M4_CDNS_5 $T=62760 161760 0 0 $X=62680 $Y=161510
X59 103 M5_M4_CDNS_5 $T=62760 167690 0 0 $X=62680 $Y=167440
X60 89 M5_M4_CDNS_5 $T=62760 169120 0 0 $X=62680 $Y=168870
X61 92 M5_M4_CDNS_5 $T=62760 175080 0 0 $X=62680 $Y=174830
X62 104 M5_M4_CDNS_5 $T=62760 234970 0 0 $X=62680 $Y=234720
X63 105 M5_M4_CDNS_5 $T=62760 240900 0 0 $X=62680 $Y=240650
X64 90 M5_M4_CDNS_5 $T=62760 242330 0 0 $X=62680 $Y=242080
X65 93 M5_M4_CDNS_5 $T=62760 248290 0 0 $X=62680 $Y=248040
X66 94 M5_M4_CDNS_5 $T=62770 81230 0 0 $X=62690 $Y=80980
X67 95 M5_M4_CDNS_5 $T=62770 154450 0 0 $X=62690 $Y=154200
X68 96 M5_M4_CDNS_5 $T=62770 227660 0 0 $X=62690 $Y=227410
X69 100 M5_M4_CDNS_5 $T=63490 16670 0 0 $X=63410 $Y=16420
X70 102 M5_M4_CDNS_5 $T=63490 89890 0 0 $X=63410 $Y=89640
X71 104 M5_M4_CDNS_5 $T=63490 163100 0 0 $X=63410 $Y=162850
X72 97 M5_M4_CDNS_5 $T=63820 12690 0 0 $X=63740 $Y=12440
X73 98 M5_M4_CDNS_5 $T=63820 85910 0 0 $X=63740 $Y=85660
X74 99 M5_M4_CDNS_5 $T=63820 159120 0 0 $X=63740 $Y=158870
X75 87 M4_M3_CDNS_6 $T=62210 216190 0 90 $X=61960 $Y=216110
X76 86 M4_M3_CDNS_6 $T=62240 142980 0 90 $X=61990 $Y=142900
X77 85 M4_M3_CDNS_6 $T=62300 69760 0 90 $X=62050 $Y=69680
X78 106 M4_M3_CDNS_6 $T=62650 125410 0 0 $X=62570 $Y=125160
X79 107 M4_M3_CDNS_6 $T=62650 198630 0 0 $X=62570 $Y=198380
X80 85 M4_M3_CDNS_6 $T=62740 103290 0 0 $X=62660 $Y=103040
X81 86 M4_M3_CDNS_6 $T=62740 176510 0 0 $X=62660 $Y=176260
X82 87 M4_M3_CDNS_6 $T=62740 249720 0 0 $X=62660 $Y=249470
X83 108 M4_M3_CDNS_6 $T=62740 271840 0 0 $X=62660 $Y=271590
X84 97 M4_M3_CDNS_6 $T=62750 87190 0 0 $X=62670 $Y=86940
X85 109 M4_M3_CDNS_6 $T=62750 111060 0 0 $X=62670 $Y=110810
X86 98 M4_M3_CDNS_6 $T=62750 160410 0 0 $X=62670 $Y=160160
X87 110 M4_M3_CDNS_6 $T=62750 184280 0 0 $X=62670 $Y=184030
X88 99 M4_M3_CDNS_6 $T=62750 233620 0 0 $X=62670 $Y=233370
X89 111 M4_M3_CDNS_6 $T=62750 257490 0 0 $X=62670 $Y=257240
X90 100 M4_M3_CDNS_6 $T=62760 88540 0 0 $X=62680 $Y=88290
X91 101 M4_M3_CDNS_6 $T=62760 94470 0 0 $X=62680 $Y=94220
X92 88 M4_M3_CDNS_6 $T=62760 95900 0 0 $X=62680 $Y=95650
X93 91 M4_M3_CDNS_6 $T=62760 101860 0 0 $X=62680 $Y=101610
X94 112 M4_M3_CDNS_6 $T=62760 118220 0 0 $X=62680 $Y=117970
X95 102 M4_M3_CDNS_6 $T=62760 161760 0 0 $X=62680 $Y=161510
X96 103 M4_M3_CDNS_6 $T=62760 167690 0 0 $X=62680 $Y=167440
X97 89 M4_M3_CDNS_6 $T=62760 169120 0 0 $X=62680 $Y=168870
X98 92 M4_M3_CDNS_6 $T=62760 175080 0 0 $X=62680 $Y=174830
X99 113 M4_M3_CDNS_6 $T=62760 191440 0 0 $X=62680 $Y=191190
X100 104 M4_M3_CDNS_6 $T=62760 234970 0 0 $X=62680 $Y=234720
X101 105 M4_M3_CDNS_6 $T=62760 240900 0 0 $X=62680 $Y=240650
X102 90 M4_M3_CDNS_6 $T=62760 242330 0 0 $X=62680 $Y=242080
X103 93 M4_M3_CDNS_6 $T=62760 248290 0 0 $X=62680 $Y=248040
X104 114 M4_M3_CDNS_6 $T=62760 264650 0 0 $X=62680 $Y=264400
X105 94 M4_M3_CDNS_6 $T=62770 81230 0 0 $X=62690 $Y=80980
X106 95 M4_M3_CDNS_6 $T=62770 154450 0 0 $X=62690 $Y=154200
X107 96 M4_M3_CDNS_6 $T=62770 227660 0 0 $X=62690 $Y=227410
X108 100 M4_M3_CDNS_6 $T=63490 16670 0 0 $X=63410 $Y=16420
X109 102 M4_M3_CDNS_6 $T=63490 89890 0 0 $X=63410 $Y=89640
X110 104 M4_M3_CDNS_6 $T=63490 163100 0 0 $X=63410 $Y=162850
X111 97 M4_M3_CDNS_6 $T=63820 12690 0 0 $X=63740 $Y=12440
X112 98 M4_M3_CDNS_6 $T=63820 85910 0 0 $X=63740 $Y=85660
X113 99 M4_M3_CDNS_6 $T=63820 159120 0 0 $X=63740 $Y=158870
X114 87 M3_M2_CDNS_7 $T=62210 216190 0 90 $X=61960 $Y=216110
X115 86 M3_M2_CDNS_7 $T=62240 142980 0 90 $X=61990 $Y=142900
X116 85 M3_M2_CDNS_7 $T=62300 69760 0 90 $X=62050 $Y=69680
X117 106 M3_M2_CDNS_7 $T=62650 125410 0 0 $X=62570 $Y=125160
X118 107 M3_M2_CDNS_7 $T=62650 198630 0 0 $X=62570 $Y=198380
X119 85 M3_M2_CDNS_7 $T=62740 103290 0 0 $X=62660 $Y=103040
X120 86 M3_M2_CDNS_7 $T=62740 176510 0 0 $X=62660 $Y=176260
X121 87 M3_M2_CDNS_7 $T=62740 249720 0 0 $X=62660 $Y=249470
X122 108 M3_M2_CDNS_7 $T=62740 271840 0 0 $X=62660 $Y=271590
X123 97 M3_M2_CDNS_7 $T=62750 87190 0 0 $X=62670 $Y=86940
X124 109 M3_M2_CDNS_7 $T=62750 111060 0 0 $X=62670 $Y=110810
X125 98 M3_M2_CDNS_7 $T=62750 160410 0 0 $X=62670 $Y=160160
X126 110 M3_M2_CDNS_7 $T=62750 184280 0 0 $X=62670 $Y=184030
X127 99 M3_M2_CDNS_7 $T=62750 233620 0 0 $X=62670 $Y=233370
X128 111 M3_M2_CDNS_7 $T=62750 257490 0 0 $X=62670 $Y=257240
X129 100 M3_M2_CDNS_7 $T=62760 88540 0 0 $X=62680 $Y=88290
X130 101 M3_M2_CDNS_7 $T=62760 94470 0 0 $X=62680 $Y=94220
X131 88 M3_M2_CDNS_7 $T=62760 95900 0 0 $X=62680 $Y=95650
X132 91 M3_M2_CDNS_7 $T=62760 101860 0 0 $X=62680 $Y=101610
X133 112 M3_M2_CDNS_7 $T=62760 118220 0 0 $X=62680 $Y=117970
X134 102 M3_M2_CDNS_7 $T=62760 161760 0 0 $X=62680 $Y=161510
X135 103 M3_M2_CDNS_7 $T=62760 167690 0 0 $X=62680 $Y=167440
X136 89 M3_M2_CDNS_7 $T=62760 169120 0 0 $X=62680 $Y=168870
X137 92 M3_M2_CDNS_7 $T=62760 175080 0 0 $X=62680 $Y=174830
X138 113 M3_M2_CDNS_7 $T=62760 191440 0 0 $X=62680 $Y=191190
X139 104 M3_M2_CDNS_7 $T=62760 234970 0 0 $X=62680 $Y=234720
X140 105 M3_M2_CDNS_7 $T=62760 240900 0 0 $X=62680 $Y=240650
X141 90 M3_M2_CDNS_7 $T=62760 242330 0 0 $X=62680 $Y=242080
X142 93 M3_M2_CDNS_7 $T=62760 248290 0 0 $X=62680 $Y=248040
X143 114 M3_M2_CDNS_7 $T=62760 264650 0 0 $X=62680 $Y=264400
X144 94 M3_M2_CDNS_7 $T=62770 81230 0 0 $X=62690 $Y=80980
X145 95 M3_M2_CDNS_7 $T=62770 154450 0 0 $X=62690 $Y=154200
X146 96 M3_M2_CDNS_7 $T=62770 227660 0 0 $X=62690 $Y=227410
X147 100 M3_M2_CDNS_7 $T=63490 16670 0 0 $X=63410 $Y=16420
X148 102 M3_M2_CDNS_7 $T=63490 89890 0 0 $X=63410 $Y=89640
X149 104 M3_M2_CDNS_7 $T=63490 163100 0 0 $X=63410 $Y=162850
X150 97 M3_M2_CDNS_7 $T=63820 12690 0 0 $X=63740 $Y=12440
X151 98 M3_M2_CDNS_7 $T=63820 85910 0 0 $X=63740 $Y=85660
X152 99 M3_M2_CDNS_7 $T=63820 159120 0 0 $X=63740 $Y=158870
X153 101 M3_M2_CDNS_7 $T=63830 19990 0 0 $X=63750 $Y=19740
X154 103 M3_M2_CDNS_7 $T=63830 93210 0 0 $X=63750 $Y=92960
X155 105 M3_M2_CDNS_7 $T=63830 166420 0 0 $X=63750 $Y=166170
X156 94 M3_M2_CDNS_7 $T=63870 9350 0 0 $X=63790 $Y=9100
X157 95 M3_M2_CDNS_7 $T=63870 82570 0 0 $X=63790 $Y=82320
X158 96 M3_M2_CDNS_7 $T=63870 155780 0 0 $X=63790 $Y=155530
X159 106 M2_M1_CDNS_8 $T=63810 53250 0 0 $X=63730 $Y=53120
X160 107 M2_M1_CDNS_8 $T=63810 126470 0 0 $X=63730 $Y=126340
X161 108 M2_M1_CDNS_8 $T=63810 199680 0 0 $X=63730 $Y=199550
X162 112 M2_M1_CDNS_8 $T=63830 45950 0 0 $X=63750 $Y=45820
X163 113 M2_M1_CDNS_8 $T=63830 119170 0 0 $X=63750 $Y=119040
X164 114 M2_M1_CDNS_8 $T=63830 192380 0 0 $X=63750 $Y=192250
X165 109 M2_M1_CDNS_8 $T=63860 38630 0 0 $X=63780 $Y=38500
X166 110 M2_M1_CDNS_8 $T=63860 111850 0 0 $X=63780 $Y=111720
X167 111 M2_M1_CDNS_8 $T=63860 185060 0 0 $X=63780 $Y=184930
X168 87 M2_M1_CDNS_9 $T=62210 216190 0 90 $X=61960 $Y=216110
X169 86 M2_M1_CDNS_9 $T=62240 142980 0 90 $X=61990 $Y=142900
X170 85 M2_M1_CDNS_9 $T=62300 69760 0 90 $X=62050 $Y=69680
X171 106 M2_M1_CDNS_9 $T=62650 125410 0 0 $X=62570 $Y=125160
X172 107 M2_M1_CDNS_9 $T=62650 198630 0 0 $X=62570 $Y=198380
X173 85 M2_M1_CDNS_9 $T=62740 103290 0 0 $X=62660 $Y=103040
X174 86 M2_M1_CDNS_9 $T=62740 176510 0 0 $X=62660 $Y=176260
X175 87 M2_M1_CDNS_9 $T=62740 249720 0 0 $X=62660 $Y=249470
X176 108 M2_M1_CDNS_9 $T=62740 271840 0 0 $X=62660 $Y=271590
X177 97 M2_M1_CDNS_9 $T=62750 87190 0 0 $X=62670 $Y=86940
X178 109 M2_M1_CDNS_9 $T=62750 111060 0 0 $X=62670 $Y=110810
X179 98 M2_M1_CDNS_9 $T=62750 160410 0 0 $X=62670 $Y=160160
X180 110 M2_M1_CDNS_9 $T=62750 184280 0 0 $X=62670 $Y=184030
X181 99 M2_M1_CDNS_9 $T=62750 233620 0 0 $X=62670 $Y=233370
X182 111 M2_M1_CDNS_9 $T=62750 257490 0 0 $X=62670 $Y=257240
X183 100 M2_M1_CDNS_9 $T=62760 88540 0 0 $X=62680 $Y=88290
X184 101 M2_M1_CDNS_9 $T=62760 94470 0 0 $X=62680 $Y=94220
X185 88 M2_M1_CDNS_9 $T=62760 95900 0 0 $X=62680 $Y=95650
X186 91 M2_M1_CDNS_9 $T=62760 101860 0 0 $X=62680 $Y=101610
X187 112 M2_M1_CDNS_9 $T=62760 118220 0 0 $X=62680 $Y=117970
X188 102 M2_M1_CDNS_9 $T=62760 161760 0 0 $X=62680 $Y=161510
X189 103 M2_M1_CDNS_9 $T=62760 167690 0 0 $X=62680 $Y=167440
X190 89 M2_M1_CDNS_9 $T=62760 169120 0 0 $X=62680 $Y=168870
X191 92 M2_M1_CDNS_9 $T=62760 175080 0 0 $X=62680 $Y=174830
X192 113 M2_M1_CDNS_9 $T=62760 191440 0 0 $X=62680 $Y=191190
X193 104 M2_M1_CDNS_9 $T=62760 234970 0 0 $X=62680 $Y=234720
X194 105 M2_M1_CDNS_9 $T=62760 240900 0 0 $X=62680 $Y=240650
X195 90 M2_M1_CDNS_9 $T=62760 242330 0 0 $X=62680 $Y=242080
X196 93 M2_M1_CDNS_9 $T=62760 248290 0 0 $X=62680 $Y=248040
X197 114 M2_M1_CDNS_9 $T=62760 264650 0 0 $X=62680 $Y=264400
X198 94 M2_M1_CDNS_9 $T=62770 81230 0 0 $X=62690 $Y=80980
X199 95 M2_M1_CDNS_9 $T=62770 154450 0 0 $X=62690 $Y=154200
X200 96 M2_M1_CDNS_9 $T=62770 227660 0 0 $X=62690 $Y=227410
X201 100 M2_M1_CDNS_9 $T=63490 16670 0 0 $X=63410 $Y=16420
X202 102 M2_M1_CDNS_9 $T=63490 89890 0 0 $X=63410 $Y=89640
X203 104 M2_M1_CDNS_9 $T=63490 163100 0 0 $X=63410 $Y=162850
X204 97 M2_M1_CDNS_9 $T=63820 12690 0 0 $X=63740 $Y=12440
X205 98 M2_M1_CDNS_9 $T=63820 85910 0 0 $X=63740 $Y=85660
X206 99 M2_M1_CDNS_9 $T=63820 159120 0 0 $X=63740 $Y=158870
X207 101 M2_M1_CDNS_9 $T=63830 19990 0 0 $X=63750 $Y=19740
X208 103 M2_M1_CDNS_9 $T=63830 93210 0 0 $X=63750 $Y=92960
X209 105 M2_M1_CDNS_9 $T=63830 166420 0 0 $X=63750 $Y=166170
X210 94 M2_M1_CDNS_9 $T=63870 9350 0 0 $X=63790 $Y=9100
X211 95 M2_M1_CDNS_9 $T=63870 82570 0 0 $X=63790 $Y=82320
X212 96 M2_M1_CDNS_9 $T=63870 155780 0 0 $X=63790 $Y=155530
X213 115 M5_M4_CDNS_10 $T=9410 93400 0 0 $X=9330 $Y=93270
X214 116 M5_M4_CDNS_10 $T=9410 166620 0 0 $X=9330 $Y=166490
X215 117 M5_M4_CDNS_10 $T=9410 239830 0 0 $X=9330 $Y=239700
X216 118 M5_M4_CDNS_10 $T=9820 94000 0 0 $X=9740 $Y=93870
X217 119 M5_M4_CDNS_10 $T=9820 167220 0 0 $X=9740 $Y=167090
X218 120 M5_M4_CDNS_10 $T=9820 240430 0 0 $X=9740 $Y=240300
X219 121 M5_M4_CDNS_10 $T=25120 73790 0 0 $X=25040 $Y=73660
X220 122 M5_M4_CDNS_10 $T=25120 147010 0 0 $X=25040 $Y=146880
X221 123 M5_M4_CDNS_10 $T=25120 220220 0 0 $X=25040 $Y=220090
X222 124 M5_M4_CDNS_10 $T=28450 130040 0 0 $X=28370 $Y=129910
X223 125 M5_M4_CDNS_10 $T=28450 203260 0 0 $X=28370 $Y=203130
X224 126 M5_M4_CDNS_10 $T=28450 276470 0 0 $X=28370 $Y=276340
X225 121 M5_M4_CDNS_10 $T=30670 73840 0 0 $X=30590 $Y=73710
X226 122 M5_M4_CDNS_10 $T=30670 147060 0 0 $X=30590 $Y=146930
X227 123 M5_M4_CDNS_10 $T=30670 220270 0 0 $X=30590 $Y=220140
X228 121 M5_M4_CDNS_10 $T=35390 130710 0 0 $X=35310 $Y=130580
X229 122 M5_M4_CDNS_10 $T=35390 203930 0 0 $X=35310 $Y=203800
X230 123 M5_M4_CDNS_10 $T=35390 277140 0 0 $X=35310 $Y=277010
X231 94 M5_M4_CDNS_10 $T=55470 70970 0 90 $X=55340 $Y=70890
X232 95 M5_M4_CDNS_10 $T=55470 144190 0 90 $X=55340 $Y=144110
X233 96 M5_M4_CDNS_10 $T=55470 217400 0 90 $X=55340 $Y=217320
X234 91 M5_M4_CDNS_10 $T=56490 100610 0 90 $X=56360 $Y=100530
X235 92 M5_M4_CDNS_10 $T=56490 173830 0 90 $X=56360 $Y=173750
X236 93 M5_M4_CDNS_10 $T=56490 247040 0 90 $X=56360 $Y=246960
X237 88 M5_M4_CDNS_10 $T=56560 97140 0 0 $X=56480 $Y=97010
X238 89 M5_M4_CDNS_10 $T=56560 170360 0 0 $X=56480 $Y=170230
X239 90 M5_M4_CDNS_10 $T=56560 243570 0 0 $X=56480 $Y=243440
X240 101 M5_M4_CDNS_10 $T=57090 92750 0 0 $X=57010 $Y=92620
X241 103 M5_M4_CDNS_10 $T=57090 165970 0 0 $X=57010 $Y=165840
X242 105 M5_M4_CDNS_10 $T=57090 239180 0 0 $X=57010 $Y=239050
X243 109 M5_M4_CDNS_10 $T=57150 110830 0 0 $X=57070 $Y=110700
X244 110 M5_M4_CDNS_10 $T=57150 184050 0 0 $X=57070 $Y=183920
X245 111 M5_M4_CDNS_10 $T=57150 257260 0 0 $X=57070 $Y=257130
X246 106 M5_M4_CDNS_10 $T=57170 125430 0 0 $X=57090 $Y=125300
X247 107 M5_M4_CDNS_10 $T=57170 198650 0 0 $X=57090 $Y=198520
X248 108 M5_M4_CDNS_10 $T=57170 271860 0 0 $X=57090 $Y=271730
X249 112 M5_M4_CDNS_10 $T=57200 118260 0 0 $X=57120 $Y=118130
X250 113 M5_M4_CDNS_10 $T=57200 191480 0 0 $X=57120 $Y=191350
X251 114 M5_M4_CDNS_10 $T=57200 264690 0 0 $X=57120 $Y=264560
X252 85 M5_M4_CDNS_10 $T=57550 103260 0 0 $X=57470 $Y=103130
X253 86 M5_M4_CDNS_10 $T=57550 176480 0 0 $X=57470 $Y=176350
X254 87 M5_M4_CDNS_10 $T=57550 249690 0 0 $X=57470 $Y=249560
X255 87 M5_M4_CDNS_10 $T=62210 216190 0 90 $X=62080 $Y=216110
X256 86 M5_M4_CDNS_10 $T=62240 142980 0 90 $X=62110 $Y=142900
X257 85 M5_M4_CDNS_10 $T=62300 69760 0 90 $X=62170 $Y=69680
X258 106 M5_M4_CDNS_10 $T=62650 125410 0 0 $X=62570 $Y=125280
X259 107 M5_M4_CDNS_10 $T=62650 198630 0 0 $X=62570 $Y=198500
X260 108 M5_M4_CDNS_10 $T=62740 271840 0 0 $X=62660 $Y=271710
X261 109 M5_M4_CDNS_10 $T=62750 111060 0 0 $X=62670 $Y=110930
X262 110 M5_M4_CDNS_10 $T=62750 184280 0 0 $X=62670 $Y=184150
X263 111 M5_M4_CDNS_10 $T=62750 257490 0 0 $X=62670 $Y=257360
X264 112 M5_M4_CDNS_10 $T=62760 118220 0 0 $X=62680 $Y=118090
X265 113 M5_M4_CDNS_10 $T=62760 191440 0 0 $X=62680 $Y=191310
X266 114 M5_M4_CDNS_10 $T=62760 264650 0 0 $X=62680 $Y=264520
X267 115 M3_M2_CDNS_11 $T=11150 139470 0 90 $X=10900 $Y=139390
X268 116 M3_M2_CDNS_11 $T=11150 212690 0 90 $X=10900 $Y=212610
X269 117 M3_M2_CDNS_11 $T=11150 285900 0 90 $X=10900 $Y=285820
X270 118 M3_M2_CDNS_11 $T=16950 140010 0 0 $X=16870 $Y=139760
X271 119 M3_M2_CDNS_11 $T=16950 213230 0 0 $X=16870 $Y=212980
X272 120 M3_M2_CDNS_11 $T=16950 286440 0 0 $X=16870 $Y=286190
X273 124 M3_M2_CDNS_11 $T=31680 139470 0 90 $X=31430 $Y=139390
X274 125 M3_M2_CDNS_11 $T=31680 212690 0 90 $X=31430 $Y=212610
X275 126 M3_M2_CDNS_11 $T=31680 285900 0 90 $X=31430 $Y=285820
X276 121 M3_M2_CDNS_11 $T=41970 139470 0 90 $X=41720 $Y=139390
X277 122 M3_M2_CDNS_11 $T=41970 212690 0 90 $X=41720 $Y=212610
X278 123 M3_M2_CDNS_11 $T=41970 285900 0 90 $X=41720 $Y=285820
X279 109 M3_M2_CDNS_11 $T=51030 71710 0 0 $X=50950 $Y=71460
X280 110 M3_M2_CDNS_11 $T=51030 144930 0 0 $X=50950 $Y=144680
X281 111 M3_M2_CDNS_11 $T=51030 218140 0 0 $X=50950 $Y=217890
X282 112 M3_M2_CDNS_11 $T=51420 72540 0 0 $X=51340 $Y=72290
X283 113 M3_M2_CDNS_11 $T=51420 145760 0 0 $X=51340 $Y=145510
X284 114 M3_M2_CDNS_11 $T=51420 218970 0 0 $X=51340 $Y=218720
X285 106 M3_M2_CDNS_11 $T=54350 80260 0 0 $X=54270 $Y=80010
X286 107 M3_M2_CDNS_11 $T=54350 153480 0 0 $X=54270 $Y=153230
X287 108 M3_M2_CDNS_11 $T=54350 226690 0 0 $X=54270 $Y=226440
X288 115 M4_M3_CDNS_12 $T=11150 139470 0 90 $X=10900 $Y=139390
X289 116 M4_M3_CDNS_12 $T=11150 212690 0 90 $X=10900 $Y=212610
X290 117 M4_M3_CDNS_12 $T=11150 285900 0 90 $X=10900 $Y=285820
X291 118 M4_M3_CDNS_12 $T=16950 140010 0 0 $X=16870 $Y=139760
X292 119 M4_M3_CDNS_12 $T=16950 213230 0 0 $X=16870 $Y=212980
X293 120 M4_M3_CDNS_12 $T=16950 286440 0 0 $X=16870 $Y=286190
X294 124 M4_M3_CDNS_12 $T=31680 139470 0 90 $X=31430 $Y=139390
X295 125 M4_M3_CDNS_12 $T=31680 212690 0 90 $X=31430 $Y=212610
X296 126 M4_M3_CDNS_12 $T=31680 285900 0 90 $X=31430 $Y=285820
X297 121 M4_M3_CDNS_12 $T=41970 139470 0 90 $X=41720 $Y=139390
X298 122 M4_M3_CDNS_12 $T=41970 212690 0 90 $X=41720 $Y=212610
X299 123 M4_M3_CDNS_12 $T=41970 285900 0 90 $X=41720 $Y=285820
X300 109 M4_M3_CDNS_12 $T=51030 71710 0 0 $X=50950 $Y=71460
X301 110 M4_M3_CDNS_12 $T=51030 144930 0 0 $X=50950 $Y=144680
X302 111 M4_M3_CDNS_12 $T=51030 218140 0 0 $X=50950 $Y=217890
X303 112 M4_M3_CDNS_12 $T=51420 72540 0 0 $X=51340 $Y=72290
X304 113 M4_M3_CDNS_12 $T=51420 145760 0 0 $X=51340 $Y=145510
X305 114 M4_M3_CDNS_12 $T=51420 218970 0 0 $X=51340 $Y=218720
X306 106 M4_M3_CDNS_12 $T=54350 80260 0 0 $X=54270 $Y=80010
X307 107 M4_M3_CDNS_12 $T=54350 153480 0 0 $X=54270 $Y=153230
X308 108 M4_M3_CDNS_12 $T=54350 226690 0 0 $X=54270 $Y=226440
X309 101 M4_M3_CDNS_12 $T=63830 19990 0 0 $X=63750 $Y=19740
X310 103 M4_M3_CDNS_12 $T=63830 93210 0 0 $X=63750 $Y=92960
X311 105 M4_M3_CDNS_12 $T=63830 166420 0 0 $X=63750 $Y=166170
X312 91 M4_M3_CDNS_13 $T=50440 71360 0 0 $X=50360 $Y=71230
X313 92 M4_M3_CDNS_13 $T=50440 144580 0 0 $X=50360 $Y=144450
X314 93 M4_M3_CDNS_13 $T=50440 217790 0 0 $X=50360 $Y=217660
X315 88 M4_M3_CDNS_13 $T=50730 70270 0 90 $X=50600 $Y=70190
X316 89 M4_M3_CDNS_13 $T=50730 143490 0 90 $X=50600 $Y=143410
X317 90 M4_M3_CDNS_13 $T=50730 216700 0 90 $X=50600 $Y=216620
X318 85 M4_M3_CDNS_13 $T=57550 91880 0 0 $X=57470 $Y=91750
X319 86 M4_M3_CDNS_13 $T=57550 165100 0 0 $X=57470 $Y=164970
X320 87 M4_M3_CDNS_13 $T=57550 238310 0 0 $X=57470 $Y=238180
X321 94 M4_M3_CDNS_13 $T=63870 9350 0 0 $X=63790 $Y=9220
X322 95 M4_M3_CDNS_13 $T=63870 82570 0 0 $X=63790 $Y=82440
X323 96 M4_M3_CDNS_13 $T=63870 155780 0 0 $X=63790 $Y=155650
X324 1 115 124 121 7 11 10 9 12 13
+ 118 8 5 6 30 36 34 35 48 43
+ 47 53 52 57 64 100 106 85 97 112
+ 101 88 109 94 91 74 73 72 71 70
+ 69 68 67 66 65 1351 2425 1271 1273 1350
+ 1347 2424 1349 1272 1314 1274 1315 1276 2423 2428
+ 1277 2427 1232 2362 1275 2430 2426 1278 1377 2466
+ 2429 1348 1346 2502 2663 2599 2600 2601 2602 2666
+ 1244 1256 1291 1302 1306 1316 1353 1354 1397 1402
+ 1420 1425 1431 1459 1477 1478 2668 2603 2604 2605
+ 2606 2670 2671 2607 2608 2609 2610 2674 2676 2611
+ 2612 2613 2614 2678 2665 2669 2673 2677 2664 2667
+ 2672 2675 ph2p2_processing_element $T=370 -60 0 0 $X=260 $Y=-60
X325 2 116 125 122 7 11 10 16 17 13
+ 119 15 115 14 31 38 118 37 49 124
+ 46 54 121 58 63 102 107 86 98 113
+ 103 89 110 95 92 94 97 100 101 88
+ 91 85 109 112 106 986 2184 906 908 985
+ 982 2183 984 907 949 909 950 911 2182 2187
+ 912 2186 867 2121 910 2189 2185 913 1012 2225
+ 2188 983 981 2261 2647 2583 2584 2585 2586 2650
+ 879 891 926 937 941 951 988 989 1032 1037
+ 1055 1060 1066 1094 1112 1113 2652 2587 2588 2589
+ 2590 2654 2655 2591 2592 2593 2594 2658 2660 2595
+ 2596 2597 2598 2662 2649 2653 2657 2661 2648 2651
+ 2656 2659 ph2p2_processing_element $T=370 73140 0 0 $X=260 $Y=73140
X326 3 117 126 123 7 11 10 20 21 13
+ 120 19 116 18 32 40 119 39 50 125
+ 45 55 122 59 62 104 108 87 99 114
+ 105 90 111 96 93 95 98 102 103 89
+ 92 86 110 113 107 621 1943 541 543 620
+ 617 1942 619 542 584 544 585 546 1941 1946
+ 547 1945 502 1880 545 1948 1944 548 647 1984
+ 1947 618 616 2020 2631 2567 2568 2569 2570 2634
+ 514 526 561 572 576 586 623 624 667 672
+ 690 695 701 729 747 748 2636 2571 2572 2573
+ 2574 2638 2639 2575 2576 2577 2578 2642 2644 2579
+ 2580 2581 2582 2646 2633 2637 2641 2645 2632 2635
+ 2640 2643 ph2p2_processing_element $T=370 146340 0 0 $X=260 $Y=146340
X327 4 25 26 27 7 11 10 28 29 13
+ 23 24 117 22 33 42 120 41 51 126
+ 44 56 123 60 61 83 75 79 77 78
+ 82 81 76 84 80 96 99 104 105 90
+ 93 87 111 114 108 256 1702 176 178 255
+ 252 1701 254 177 219 179 220 181 1700 1705
+ 182 1704 137 1639 180 1707 1703 183 282 1743
+ 1706 253 251 1779 2615 2551 2552 2553 2554 2618
+ 149 161 196 207 211 221 258 259 302 307
+ 325 330 336 364 382 383 2620 2555 2556 2557
+ 2558 2622 2623 2559 2560 2561 2562 2626 2628 2563
+ 2564 2565 2566 2630 2617 2621 2625 2629 2616 2619
+ 2624 2627 ph2p2_processing_element $T=370 219540 0 0 $X=260 $Y=219540
M0 2602 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=72010 $dt=1
M1 2586 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=145210 $dt=1
M2 2570 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=13.1038 scb=0.0126439 scc=0.000226416 $X=2290 $Y=218410 $dt=1
M3 2554 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=15.5779 scb=0.0149308 scc=0.000240309 $X=2290 $Y=291610 $dt=1
M4 1256 1232 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.8911 scb=0.00996238 scc=0.000256798 $X=2380 $Y=920 $dt=1
M5 891 867 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=74120 $dt=1
M6 526 502 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=147320 $dt=1
M7 161 137 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.90193 scb=0.0083839 scc=0.000250634 $X=2380 $Y=220520 $dt=1
M8 2663 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=72040 $dt=1
M9 2647 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=145240 $dt=1
M10 2631 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=3620 $Y=218440 $dt=1
M11 2615 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=3620 $Y=291640 $dt=1
M12 2664 1232 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=3710 $Y=680 $dt=1
M13 2648 867 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=73880 $dt=1
M14 2632 502 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=147080 $dt=1
M15 2616 137 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=3710 $Y=220280 $dt=1
M16 1291 1244 2664 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=4680 $Y=620 $dt=1
M17 926 879 2648 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=73820 $dt=1
M18 561 514 2632 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=147020 $dt=1
M19 196 149 2616 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=4680 $Y=220220 $dt=1
M20 2599 10 115 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=72040 $dt=1
M21 2583 10 116 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=145240 $dt=1
M22 2567 10 117 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=4800 $Y=218440 $dt=1
M23 2551 10 25 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=4800 $Y=291640 $dt=1
M24 1291 1256 2664 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=5640 $Y=620 $dt=1
M25 926 891 2648 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=73820 $dt=1
M26 561 526 2632 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=147020 $dt=1
M27 196 161 2616 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=5640 $Y=220220 $dt=1
M28 2601 2599 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=71950 $dt=1
M29 2585 2583 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=145150 $dt=1
M30 2569 2567 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=6000 $Y=218350 $dt=1
M31 2553 2551 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=6000 $Y=291550 $dt=1
M32 2664 12 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=6600 $Y=620 $dt=1
M33 2648 17 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=73820 $dt=1
M34 2632 21 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=147020 $dt=1
M35 2616 29 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=6600 $Y=220220 $dt=1
M36 2601 2600 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=71960 $dt=1
M37 2585 2584 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=145160 $dt=1
M38 2569 2568 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=7240 $Y=218360 $dt=1
M39 2553 2552 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=7240 $Y=291560 $dt=1
M40 1302 1316 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=8260 $Y=920 $dt=1
M41 937 951 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=74120 $dt=1
M42 572 586 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=147320 $dt=1
M43 207 221 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=8260 $Y=220520 $dt=1
M44 2665 2601 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=72010 $dt=1
M45 2649 2585 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=145210 $dt=1
M46 2633 2569 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=8490 $Y=218410 $dt=1
M47 2617 2553 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=8490 $Y=291610 $dt=1
M48 1306 1291 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=9220 $Y=920 $dt=1
M49 941 926 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=74120 $dt=1
M50 576 561 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=147320 $dt=1
M51 211 196 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=9220 $Y=220520 $dt=1
M52 2666 2602 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=72040 $dt=1
M53 2650 2586 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=145240 $dt=1
M54 2634 2570 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=9820 $Y=218440 $dt=1
M55 2618 2554 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=9820 $Y=291640 $dt=1
M56 2667 1291 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=10550 $Y=680 $dt=1
M57 2651 926 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=73880 $dt=1
M58 2635 561 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=147080 $dt=1
M59 2619 196 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=10550 $Y=220280 $dt=1
M60 2599 2602 2665 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=72040 $dt=1
M61 2583 2586 2649 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=145240 $dt=1
M62 2567 2570 2633 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=11000 $Y=218440 $dt=1
M63 2551 2554 2617 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=11000 $Y=291640 $dt=1
M64 2362 1302 2667 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=11520 $Y=620 $dt=1
M65 2121 937 2651 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=73820 $dt=1
M66 1880 572 2635 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=147020 $dt=1
M67 1639 207 2619 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=11520 $Y=220220 $dt=1
M68 2362 1306 2667 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=12480 $Y=620 $dt=1
M69 2121 941 2651 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=73820 $dt=1
M70 1880 576 2635 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=147020 $dt=1
M71 1639 211 2619 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=12480 $Y=220220 $dt=1
M72 2606 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=72010 $dt=1
M73 2590 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=145210 $dt=1
M74 2574 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=12530 $Y=218410 $dt=1
M75 2558 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=12530 $Y=291610 $dt=1
M76 2667 1316 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=13440 $Y=620 $dt=1
M77 2651 951 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=73820 $dt=1
M78 2635 586 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=147020 $dt=1
M79 2619 221 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=13440 $Y=220220 $dt=1
M80 2668 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=72040 $dt=1
M81 2652 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=145240 $dt=1
M82 2636 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=13860 $Y=218440 $dt=1
M83 2620 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=13860 $Y=291640 $dt=1
M84 2603 10 118 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=72040 $dt=1
M85 2587 10 119 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=145240 $dt=1
M86 2571 10 120 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=15040 $Y=218440 $dt=1
M87 2555 10 23 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=15040 $Y=291640 $dt=1
M88 1353 1316 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=15510 $Y=650 $dt=1
M89 988 951 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=73850 $dt=1
M90 623 586 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=147050 $dt=1
M91 258 221 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15510 $Y=220250 $dt=1
M92 13 1291 1353 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=15920 $Y=650 $dt=1
M93 13 926 988 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=73850 $dt=1
M94 13 561 623 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=147050 $dt=1
M95 13 196 258 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=15920 $Y=220250 $dt=1
M96 2605 2603 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=71950 $dt=1
M97 2589 2587 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=145150 $dt=1
M98 2573 2571 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=16240 $Y=218350 $dt=1
M99 2557 2555 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=16240 $Y=291550 $dt=1
M100 2605 2604 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=71960 $dt=1
M101 2589 2588 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=145160 $dt=1
M102 2573 2572 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=17480 $Y=218360 $dt=1
M103 2557 2556 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=17480 $Y=291560 $dt=1
M104 1354 12 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=18490 $Y=910 $dt=1
M105 989 17 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=74110 $dt=1
M106 624 21 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=147310 $dt=1
M107 259 29 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18490 $Y=220510 $dt=1
M108 2669 2605 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=72010 $dt=1
M109 2653 2589 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=145210 $dt=1
M110 2637 2573 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=18730 $Y=218410 $dt=1
M111 2621 2557 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=18730 $Y=291610 $dt=1
M112 13 1232 1354 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=18900 $Y=910 $dt=1
M113 13 867 989 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=74110 $dt=1
M114 13 502 624 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=147310 $dt=1
M115 13 137 259 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=18900 $Y=220510 $dt=1
M116 2670 2606 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=72040 $dt=1
M117 2654 2590 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=145240 $dt=1
M118 2638 2574 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=20060 $Y=218440 $dt=1
M119 2622 2558 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=20060 $Y=291640 $dt=1
M120 2603 2606 2669 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=72040 $dt=1
M121 2587 2590 2653 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=145240 $dt=1
M122 2571 2574 2637 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=21240 $Y=218440 $dt=1
M123 2555 2558 2621 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=21240 $Y=291640 $dt=1
M124 1459 1353 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=21330 $Y=910 $dt=1
M125 1094 988 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=74110 $dt=1
M126 729 623 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=147310 $dt=1
M127 364 258 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21330 $Y=220510 $dt=1
M128 13 1354 1459 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=21740 $Y=910 $dt=1
M129 13 989 1094 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=74110 $dt=1
M130 13 624 729 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=147310 $dt=1
M131 13 259 364 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=21740 $Y=220510 $dt=1
M132 2610 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=72010 $dt=1
M133 2594 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=145210 $dt=1
M134 2578 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=22770 $Y=218410 $dt=1
M135 2562 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=22770 $Y=291610 $dt=1
M136 1397 48 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=23380 $Y=920 $dt=1
M137 1032 49 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=74120 $dt=1
M138 667 50 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=147320 $dt=1
M139 302 51 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=23380 $Y=220520 $dt=1
M140 2671 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=72040 $dt=1
M141 2655 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=145240 $dt=1
M142 2639 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=24100 $Y=218440 $dt=1
M143 2623 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=24100 $Y=291640 $dt=1
M144 1402 1377 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=24340 $Y=920 $dt=1
M145 1037 1012 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=74120 $dt=1
M146 672 647 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=147320 $dt=1
M147 307 282 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=24340 $Y=220520 $dt=1
M148 2607 10 124 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=72040 $dt=1
M149 2591 10 125 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=145240 $dt=1
M150 2575 10 126 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=25280 $Y=218440 $dt=1
M151 2559 10 26 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=25280 $Y=291640 $dt=1
M152 2672 1377 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=25670 $Y=680 $dt=1
M153 2656 1012 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=73880 $dt=1
M154 2640 647 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=147080 $dt=1
M155 2624 282 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=25670 $Y=220280 $dt=1
M156 2609 2607 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=71950 $dt=1
M157 2593 2591 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=145150 $dt=1
M158 2577 2575 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=26480 $Y=218350 $dt=1
M159 2561 2559 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=26480 $Y=291550 $dt=1
M160 1420 1397 2672 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=26640 $Y=620 $dt=1
M161 1055 1032 2656 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=73820 $dt=1
M162 690 667 2640 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=147020 $dt=1
M163 325 302 2624 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=26640 $Y=220220 $dt=1
M164 1420 1402 2672 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=27600 $Y=620 $dt=1
M165 1055 1037 2656 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=73820 $dt=1
M166 690 672 2640 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=147020 $dt=1
M167 325 307 2624 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=27600 $Y=220220 $dt=1
M168 2609 2608 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=71960 $dt=1
M169 2593 2592 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=145160 $dt=1
M170 2577 2576 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=27720 $Y=218360 $dt=1
M171 2561 2560 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=27720 $Y=291560 $dt=1
M172 2672 48 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=28560 $Y=620 $dt=1
M173 2656 49 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=73820 $dt=1
M174 2640 50 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=147020 $dt=1
M175 2624 51 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=28560 $Y=220220 $dt=1
M176 2673 2609 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=72010 $dt=1
M177 2657 2593 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=145210 $dt=1
M178 2641 2577 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=28970 $Y=218410 $dt=1
M179 2625 2561 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=28970 $Y=291610 $dt=1
M180 1425 1459 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=30220 $Y=920 $dt=1
M181 1060 1094 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=74120 $dt=1
M182 695 729 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=147320 $dt=1
M183 330 364 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=30220 $Y=220520 $dt=1
M184 2674 2610 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=72040 $dt=1
M185 2658 2594 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=145240 $dt=1
M186 2642 2578 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=30300 $Y=218440 $dt=1
M187 2626 2562 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=30300 $Y=291640 $dt=1
M188 1431 1420 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.5776 scb=0.00987478 scc=0.000256781 $X=31180 $Y=920 $dt=1
M189 1066 1055 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=74120 $dt=1
M190 701 690 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=147320 $dt=1
M191 336 325 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.58846 scb=0.0082963 scc=0.000250617 $X=31180 $Y=220520 $dt=1
M192 2607 2610 2673 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=72040 $dt=1
M193 2591 2594 2657 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=145240 $dt=1
M194 2575 2578 2641 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=31480 $Y=218440 $dt=1
M195 2559 2562 2625 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=31480 $Y=291640 $dt=1
M196 2675 1420 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=14.8592 scb=0.0131351 scc=0.000918216 $X=32510 $Y=680 $dt=1
M197 2659 1055 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=73880 $dt=1
M198 2643 690 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=147080 $dt=1
M199 2627 325 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=12.3552 scb=0.0107648 scc=0.000891478 $X=32510 $Y=220280 $dt=1
M200 2614 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=72010 $dt=1
M201 2598 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=145210 $dt=1
M202 2582 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=33010 $Y=218410 $dt=1
M203 2566 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=33010 $Y=291610 $dt=1
M204 2466 1425 2675 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=33480 $Y=620 $dt=1
M205 2225 1060 2659 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=73820 $dt=1
M206 1984 695 2643 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=147020 $dt=1
M207 1743 330 2627 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=33480 $Y=220220 $dt=1
M208 2676 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=72040 $dt=1
M209 2660 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=145240 $dt=1
M210 2644 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.79132 scb=0.00535378 scc=8.92944e-05 $X=34340 $Y=218440 $dt=1
M211 2628 10 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.4559 scb=0.00793674 scc=0.000107477 $X=34340 $Y=291640 $dt=1
M212 2466 1431 2675 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=34440 $Y=620 $dt=1
M213 2225 1066 2659 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=73820 $dt=1
M214 1984 701 2643 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=147020 $dt=1
M215 1743 336 2627 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=34440 $Y=220220 $dt=1
M216 2675 1459 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=13.3561 scb=0.0119202 scc=0.000604399 $X=35400 $Y=620 $dt=1
M217 2659 1094 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=73820 $dt=1
M218 2643 729 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=147020 $dt=1
M219 2627 364 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=6.72e-14 PD=1.24e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=1.4e-07 sca=10.445 scb=0.0089239 scc=0.000559159 $X=35400 $Y=220220 $dt=1
M220 2611 10 121 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=72040 $dt=1
M221 2595 10 122 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=145240 $dt=1
M222 2579 10 123 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=9.20059 scb=0.00764836 scc=0.000159521 $X=35520 $Y=218440 $dt=1
M223 2563 10 27 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0214 scb=0.00904448 scc=0.000163241 $X=35520 $Y=291640 $dt=1
M224 2613 2611 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=71950 $dt=1
M225 2597 2595 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=145150 $dt=1
M226 2581 2579 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=9.05646 scb=0.00745111 scc=0.000194153 $X=36720 $Y=218350 $dt=1
M227 2565 2563 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.1944 scb=0.00923888 scc=0.000202241 $X=36720 $Y=291550 $dt=1
M228 1477 1459 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=37470 $Y=650 $dt=1
M229 1112 1094 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=73850 $dt=1
M230 747 729 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=147050 $dt=1
M231 382 364 13 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=7.68e-14 AS=6.72e-14 PD=1.28e-06 PS=1.24e-06 fw=4.8e-07 sa=1.4e-07 sb=3.45e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37470 $Y=220250 $dt=1
M232 13 1420 1477 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=14.0115 scb=0.0124823 scc=0.000742408 $X=37880 $Y=650 $dt=1
M233 13 1055 1112 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=73850 $dt=1
M234 13 690 747 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=147050 $dt=1
M235 13 325 382 13 g45p1svt L=4.5e-08 W=4.8e-07 AD=6.72e-14 AS=7.68e-14 PD=1.24e-06 PS=1.28e-06 fw=4.8e-07 sa=3.45e-07 sb=1.4e-07 sca=11.3137 scb=0.00981578 scc=0.000707604 $X=37880 $Y=220250 $dt=1
M236 2613 2612 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=71960 $dt=1
M237 2597 2596 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=145160 $dt=1
M238 2581 2580 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.89317 scb=0.00718657 scc=0.000178238 $X=37960 $Y=218360 $dt=1
M239 2565 2564 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=11.0834 scb=0.00904972 scc=0.000187092 $X=37960 $Y=291560 $dt=1
M240 2677 2613 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=72010 $dt=1
M241 2661 2597 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=145210 $dt=1
M242 2645 2581 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=8.16621 scb=0.00598477 scc=0.000115874 $X=39210 $Y=218410 $dt=1
M243 2629 2565 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6403 scb=0.00827174 scc=0.000129767 $X=39210 $Y=291610 $dt=1
M244 1478 48 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=40450 $Y=910 $dt=1
M245 1113 49 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=74110 $dt=1
M246 748 50 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=147310 $dt=1
M247 383 51 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.84e-14 AS=3.36e-14 PD=8e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=3.45e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40450 $Y=220510 $dt=1
M248 2678 2614 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=72040 $dt=1
M249 2662 2598 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=145240 $dt=1
M250 2646 2582 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=7.96076 scb=0.005393 scc=8.92993e-05 $X=40540 $Y=218440 $dt=1
M251 2630 2566 13 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.36e-14 PD=7.6e-07 PS=7.6e-07 fw=2.4e-07 sa=1.4e-07 sb=1.4e-07 sca=10.6253 scb=0.00797597 scc=0.000107482 $X=40540 $Y=291640 $dt=1
M252 13 1377 1478 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=11.4412 scb=0.00965134 scc=0.000236974 $X=40860 $Y=910 $dt=1
M253 13 1012 1113 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=74110 $dt=1
M254 13 647 748 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=147310 $dt=1
M255 13 282 383 13 g45p1svt L=4.5e-08 W=2.4e-07 AD=3.36e-14 AS=3.84e-14 PD=7.6e-07 PS=8e-07 fw=2.4e-07 sa=3.45e-07 sb=1.4e-07 sca=9.4037 scb=0.0080058 scc=0.000230225 $X=40860 $Y=220510 $dt=1
M256 2611 2614 2677 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=72040 $dt=1
M257 2595 2598 2661 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=145240 $dt=1
M258 2579 2582 2645 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=16.3245 scb=0.0180307 scc=0.000472719 $X=41720 $Y=218440 $dt=1
M259 2563 2566 2629 13 g45p1svt L=4.5e-08 W=1.2e-07 AD=1.68e-14 AS=1.68e-14 PD=5.2e-07 PS=5.2e-07 fw=1.2e-07 sa=1.4e-07 sb=1.4e-07 sca=18.1453 scb=0.0194268 scc=0.000476439 $X=41720 $Y=291640 $dt=1
.ends ph2p3_Matrix_vector_Multiplication

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ph3_sytolic_array                               *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ph3_sytolic_array 94 85 99 79 78 98 89 75 97 66
+ 71 96 240 228 226 216 93 137 143 76
+ 131 142 88 129 141 65 127 140 239 229
+ 225 212 92 177 183 73 171 182 87 169
+ 181 64 167 180 238 230 224 209 91 221
+ 235 68 214 234 86 211 233 63 208 232
+ 237 231 223 206 81 80 82 83 67 90
+ 95 100 133 132 134 135 125 138 139 144
+ 173 172 174 175 165 178 179 184 217 215
+ 218 219 205 222 227 236 2 84 77 74
+ 70 136 130 128 126 176 170 168 166 220
+ 213 210 207 1 104 103 102 101 105 106
+ 107 108 110 112 114 109 111 113 115 118
+ 116 119 121 123 124 120 122 117 145 146
+ 147 148 150 152 154 149 151 153 155 158
+ 156 159 161 163 164 160 162 157 185 186
+ 187 188 190 192 194 189 191 193 195 198
+ 196 199 201 203 204 200 202 197 245 246
+ 247 248 250 252 254 249 251 253 255 258
+ 256 259 261 263 264 260 262 257 69 241
+ 242 243 244 72
** N=10128 EP=204 FDC=26592
X0 1 M3_M2_CDNS_1 $T=34030 66930 0 0 $X=33950 $Y=66680
X1 1 M3_M2_CDNS_1 $T=34030 68540 0 0 $X=33950 $Y=68290
X2 1 M3_M2_CDNS_1 $T=34030 140130 0 0 $X=33950 $Y=139880
X3 1 M3_M2_CDNS_1 $T=34030 141740 0 0 $X=33950 $Y=141490
X4 1 M3_M2_CDNS_1 $T=34030 213330 0 0 $X=33950 $Y=213080
X5 1 M3_M2_CDNS_1 $T=34030 214940 0 0 $X=33950 $Y=214690
X6 1 M3_M2_CDNS_1 $T=34030 286530 0 0 $X=33950 $Y=286280
X7 1 M3_M2_CDNS_1 $T=34030 288140 0 0 $X=33950 $Y=287890
X8 2 M3_M2_CDNS_1 $T=48420 72600 0 0 $X=48340 $Y=72350
X9 2 M3_M2_CDNS_1 $T=48420 145800 0 0 $X=48340 $Y=145550
X10 2 M3_M2_CDNS_1 $T=48420 219000 0 0 $X=48340 $Y=218750
X11 3 M3_M2_CDNS_1 $T=48580 60970 0 0 $X=48500 $Y=60720
X12 4 M3_M2_CDNS_1 $T=48580 134170 0 0 $X=48500 $Y=133920
X13 5 M3_M2_CDNS_1 $T=48580 207370 0 0 $X=48500 $Y=207120
X14 6 M3_M2_CDNS_1 $T=48610 60050 0 0 $X=48530 $Y=59800
X15 7 M3_M2_CDNS_1 $T=48610 133250 0 0 $X=48530 $Y=133000
X16 8 M3_M2_CDNS_1 $T=48610 206450 0 0 $X=48530 $Y=206200
X17 9 M3_M2_CDNS_1 $T=48640 59100 0 0 $X=48560 $Y=58850
X18 10 M3_M2_CDNS_1 $T=48640 132300 0 0 $X=48560 $Y=132050
X19 11 M3_M2_CDNS_1 $T=48640 205500 0 0 $X=48560 $Y=205250
X20 12 M3_M2_CDNS_1 $T=48710 65320 0 0 $X=48630 $Y=65070
X21 13 M3_M2_CDNS_1 $T=48710 138520 0 0 $X=48630 $Y=138270
X22 14 M3_M2_CDNS_1 $T=48710 211720 0 0 $X=48630 $Y=211470
X23 1 M3_M2_CDNS_1 $T=61670 68120 0 0 $X=61590 $Y=67870
X24 1 M3_M2_CDNS_1 $T=61670 141320 0 0 $X=61590 $Y=141070
X25 1 M3_M2_CDNS_1 $T=61670 214520 0 0 $X=61590 $Y=214270
X26 1 M3_M2_CDNS_1 $T=63700 68120 0 0 $X=63620 $Y=67870
X27 1 M3_M2_CDNS_1 $T=63700 141320 0 0 $X=63620 $Y=141070
X28 1 M3_M2_CDNS_1 $T=63700 214520 0 0 $X=63620 $Y=214270
X29 3 M3_M2_CDNS_1 $T=63840 57970 0 0 $X=63760 $Y=57720
X30 4 M3_M2_CDNS_1 $T=63840 131170 0 0 $X=63760 $Y=130920
X31 5 M3_M2_CDNS_1 $T=63840 204370 0 0 $X=63760 $Y=204120
X32 6 M3_M2_CDNS_1 $T=64280 60020 0 0 $X=64200 $Y=59770
X33 7 M3_M2_CDNS_1 $T=64280 133220 0 0 $X=64200 $Y=132970
X34 8 M3_M2_CDNS_1 $T=64280 206420 0 0 $X=64200 $Y=206170
X35 1 M3_M2_CDNS_1 $T=98120 66930 0 0 $X=98040 $Y=66680
X36 1 M3_M2_CDNS_1 $T=98120 68540 0 0 $X=98040 $Y=68290
X37 1 M3_M2_CDNS_1 $T=98120 140130 0 0 $X=98040 $Y=139880
X38 1 M3_M2_CDNS_1 $T=98120 141740 0 0 $X=98040 $Y=141490
X39 1 M3_M2_CDNS_1 $T=98120 213330 0 0 $X=98040 $Y=213080
X40 1 M3_M2_CDNS_1 $T=98120 214940 0 0 $X=98040 $Y=214690
X41 1 M3_M2_CDNS_1 $T=98120 286530 0 0 $X=98040 $Y=286280
X42 1 M3_M2_CDNS_1 $T=98120 288140 0 0 $X=98040 $Y=287890
X43 2 M3_M2_CDNS_1 $T=112510 72600 0 0 $X=112430 $Y=72350
X44 2 M3_M2_CDNS_1 $T=112510 145800 0 0 $X=112430 $Y=145550
X45 2 M3_M2_CDNS_1 $T=112510 219000 0 0 $X=112430 $Y=218750
X46 15 M3_M2_CDNS_1 $T=112670 60970 0 0 $X=112590 $Y=60720
X47 16 M3_M2_CDNS_1 $T=112670 134170 0 0 $X=112590 $Y=133920
X48 17 M3_M2_CDNS_1 $T=112670 207370 0 0 $X=112590 $Y=207120
X49 18 M3_M2_CDNS_1 $T=112700 60050 0 0 $X=112620 $Y=59800
X50 19 M3_M2_CDNS_1 $T=112700 133250 0 0 $X=112620 $Y=133000
X51 20 M3_M2_CDNS_1 $T=112700 206450 0 0 $X=112620 $Y=206200
X52 21 M3_M2_CDNS_1 $T=112730 59100 0 0 $X=112650 $Y=58850
X53 22 M3_M2_CDNS_1 $T=112730 132300 0 0 $X=112650 $Y=132050
X54 23 M3_M2_CDNS_1 $T=112730 205500 0 0 $X=112650 $Y=205250
X55 24 M3_M2_CDNS_1 $T=112800 65320 0 0 $X=112720 $Y=65070
X56 25 M3_M2_CDNS_1 $T=112800 138520 0 0 $X=112720 $Y=138270
X57 26 M3_M2_CDNS_1 $T=112800 211720 0 0 $X=112720 $Y=211470
X58 27 M3_M2_CDNS_1 $T=114770 6460 0 0 $X=114690 $Y=6210
X59 28 M3_M2_CDNS_1 $T=114770 79660 0 0 $X=114690 $Y=79410
X60 29 M3_M2_CDNS_1 $T=114770 152860 0 0 $X=114690 $Y=152610
X61 30 M3_M2_CDNS_1 $T=114770 226060 0 0 $X=114690 $Y=225810
X62 1 M3_M2_CDNS_1 $T=125760 68120 0 0 $X=125680 $Y=67870
X63 1 M3_M2_CDNS_1 $T=125760 141320 0 0 $X=125680 $Y=141070
X64 1 M3_M2_CDNS_1 $T=125760 214520 0 0 $X=125680 $Y=214270
X65 1 M3_M2_CDNS_1 $T=127790 68120 0 0 $X=127710 $Y=67870
X66 1 M3_M2_CDNS_1 $T=127790 141320 0 0 $X=127710 $Y=141070
X67 1 M3_M2_CDNS_1 $T=127790 214520 0 0 $X=127710 $Y=214270
X68 15 M3_M2_CDNS_1 $T=127930 57970 0 0 $X=127850 $Y=57720
X69 16 M3_M2_CDNS_1 $T=127930 131170 0 0 $X=127850 $Y=130920
X70 17 M3_M2_CDNS_1 $T=127930 204370 0 0 $X=127850 $Y=204120
X71 18 M3_M2_CDNS_1 $T=128370 60020 0 0 $X=128290 $Y=59770
X72 19 M3_M2_CDNS_1 $T=128370 133220 0 0 $X=128290 $Y=132970
X73 20 M3_M2_CDNS_1 $T=128370 206420 0 0 $X=128290 $Y=206170
X74 1 M3_M2_CDNS_1 $T=162210 66930 0 0 $X=162130 $Y=66680
X75 1 M3_M2_CDNS_1 $T=162210 68540 0 0 $X=162130 $Y=68290
X76 1 M3_M2_CDNS_1 $T=162210 140130 0 0 $X=162130 $Y=139880
X77 1 M3_M2_CDNS_1 $T=162210 141740 0 0 $X=162130 $Y=141490
X78 1 M3_M2_CDNS_1 $T=162210 213330 0 0 $X=162130 $Y=213080
X79 1 M3_M2_CDNS_1 $T=162210 214940 0 0 $X=162130 $Y=214690
X80 1 M3_M2_CDNS_1 $T=162210 286530 0 0 $X=162130 $Y=286280
X81 1 M3_M2_CDNS_1 $T=162210 288140 0 0 $X=162130 $Y=287890
X82 2 M3_M2_CDNS_1 $T=176600 72600 0 0 $X=176520 $Y=72350
X83 2 M3_M2_CDNS_1 $T=176600 145800 0 0 $X=176520 $Y=145550
X84 2 M3_M2_CDNS_1 $T=176600 219000 0 0 $X=176520 $Y=218750
X85 31 M3_M2_CDNS_1 $T=176760 60970 0 0 $X=176680 $Y=60720
X86 32 M3_M2_CDNS_1 $T=176760 134170 0 0 $X=176680 $Y=133920
X87 33 M3_M2_CDNS_1 $T=176760 207370 0 0 $X=176680 $Y=207120
X88 34 M3_M2_CDNS_1 $T=176790 60050 0 0 $X=176710 $Y=59800
X89 35 M3_M2_CDNS_1 $T=176790 133250 0 0 $X=176710 $Y=133000
X90 36 M3_M2_CDNS_1 $T=176790 206450 0 0 $X=176710 $Y=206200
X91 37 M3_M2_CDNS_1 $T=176820 59100 0 0 $X=176740 $Y=58850
X92 38 M3_M2_CDNS_1 $T=176820 132300 0 0 $X=176740 $Y=132050
X93 39 M3_M2_CDNS_1 $T=176820 205500 0 0 $X=176740 $Y=205250
X94 40 M3_M2_CDNS_1 $T=176890 65320 0 0 $X=176810 $Y=65070
X95 41 M3_M2_CDNS_1 $T=176890 138520 0 0 $X=176810 $Y=138270
X96 42 M3_M2_CDNS_1 $T=176890 211720 0 0 $X=176810 $Y=211470
X97 43 M3_M2_CDNS_1 $T=178860 6460 0 0 $X=178780 $Y=6210
X98 44 M3_M2_CDNS_1 $T=178860 79660 0 0 $X=178780 $Y=79410
X99 45 M3_M2_CDNS_1 $T=178860 152860 0 0 $X=178780 $Y=152610
X100 46 M3_M2_CDNS_1 $T=178860 226060 0 0 $X=178780 $Y=225810
X101 1 M3_M2_CDNS_1 $T=189850 68120 0 0 $X=189770 $Y=67870
X102 1 M3_M2_CDNS_1 $T=189850 141320 0 0 $X=189770 $Y=141070
X103 1 M3_M2_CDNS_1 $T=189850 214520 0 0 $X=189770 $Y=214270
X104 1 M3_M2_CDNS_1 $T=191880 68120 0 0 $X=191800 $Y=67870
X105 1 M3_M2_CDNS_1 $T=191880 141320 0 0 $X=191800 $Y=141070
X106 1 M3_M2_CDNS_1 $T=191880 214520 0 0 $X=191800 $Y=214270
X107 31 M3_M2_CDNS_1 $T=192020 57970 0 0 $X=191940 $Y=57720
X108 32 M3_M2_CDNS_1 $T=192020 131170 0 0 $X=191940 $Y=130920
X109 33 M3_M2_CDNS_1 $T=192020 204370 0 0 $X=191940 $Y=204120
X110 34 M3_M2_CDNS_1 $T=192460 60020 0 0 $X=192380 $Y=59770
X111 35 M3_M2_CDNS_1 $T=192460 133220 0 0 $X=192380 $Y=132970
X112 36 M3_M2_CDNS_1 $T=192460 206420 0 0 $X=192380 $Y=206170
X113 47 M3_M2_CDNS_1 $T=242950 6460 0 0 $X=242870 $Y=6210
X114 48 M3_M2_CDNS_1 $T=242950 79660 0 0 $X=242870 $Y=79410
X115 49 M3_M2_CDNS_1 $T=242950 152860 0 0 $X=242870 $Y=152610
X116 50 M3_M2_CDNS_1 $T=242950 226060 0 0 $X=242870 $Y=225810
X117 1 M2_M1_CDNS_2 $T=34030 66930 0 0 $X=33950 $Y=66680
X118 1 M2_M1_CDNS_2 $T=34030 68540 0 0 $X=33950 $Y=68290
X119 1 M2_M1_CDNS_2 $T=34030 140130 0 0 $X=33950 $Y=139880
X120 1 M2_M1_CDNS_2 $T=34030 141740 0 0 $X=33950 $Y=141490
X121 1 M2_M1_CDNS_2 $T=34030 213330 0 0 $X=33950 $Y=213080
X122 1 M2_M1_CDNS_2 $T=34030 214940 0 0 $X=33950 $Y=214690
X123 1 M2_M1_CDNS_2 $T=34030 286530 0 0 $X=33950 $Y=286280
X124 1 M2_M1_CDNS_2 $T=34030 288140 0 0 $X=33950 $Y=287890
X125 2 M2_M1_CDNS_2 $T=48420 72600 0 0 $X=48340 $Y=72350
X126 2 M2_M1_CDNS_2 $T=48420 145800 0 0 $X=48340 $Y=145550
X127 2 M2_M1_CDNS_2 $T=48420 219000 0 0 $X=48340 $Y=218750
X128 3 M2_M1_CDNS_2 $T=48580 60970 0 0 $X=48500 $Y=60720
X129 4 M2_M1_CDNS_2 $T=48580 134170 0 0 $X=48500 $Y=133920
X130 5 M2_M1_CDNS_2 $T=48580 207370 0 0 $X=48500 $Y=207120
X131 6 M2_M1_CDNS_2 $T=48610 60050 0 0 $X=48530 $Y=59800
X132 7 M2_M1_CDNS_2 $T=48610 133250 0 0 $X=48530 $Y=133000
X133 8 M2_M1_CDNS_2 $T=48610 206450 0 0 $X=48530 $Y=206200
X134 9 M2_M1_CDNS_2 $T=48640 59100 0 0 $X=48560 $Y=58850
X135 10 M2_M1_CDNS_2 $T=48640 132300 0 0 $X=48560 $Y=132050
X136 11 M2_M1_CDNS_2 $T=48640 205500 0 0 $X=48560 $Y=205250
X137 12 M2_M1_CDNS_2 $T=48710 65320 0 0 $X=48630 $Y=65070
X138 13 M2_M1_CDNS_2 $T=48710 138520 0 0 $X=48630 $Y=138270
X139 14 M2_M1_CDNS_2 $T=48710 211720 0 0 $X=48630 $Y=211470
X140 1 M2_M1_CDNS_2 $T=61670 68120 0 0 $X=61590 $Y=67870
X141 1 M2_M1_CDNS_2 $T=61670 141320 0 0 $X=61590 $Y=141070
X142 1 M2_M1_CDNS_2 $T=61670 214520 0 0 $X=61590 $Y=214270
X143 1 M2_M1_CDNS_2 $T=63700 68120 0 0 $X=63620 $Y=67870
X144 1 M2_M1_CDNS_2 $T=63700 141320 0 0 $X=63620 $Y=141070
X145 1 M2_M1_CDNS_2 $T=63700 214520 0 0 $X=63620 $Y=214270
X146 3 M2_M1_CDNS_2 $T=63840 57970 0 0 $X=63760 $Y=57720
X147 4 M2_M1_CDNS_2 $T=63840 131170 0 0 $X=63760 $Y=130920
X148 5 M2_M1_CDNS_2 $T=63840 204370 0 0 $X=63760 $Y=204120
X149 6 M2_M1_CDNS_2 $T=64280 60020 0 0 $X=64200 $Y=59770
X150 7 M2_M1_CDNS_2 $T=64280 133220 0 0 $X=64200 $Y=132970
X151 8 M2_M1_CDNS_2 $T=64280 206420 0 0 $X=64200 $Y=206170
X152 1 M2_M1_CDNS_2 $T=98120 66930 0 0 $X=98040 $Y=66680
X153 1 M2_M1_CDNS_2 $T=98120 68540 0 0 $X=98040 $Y=68290
X154 1 M2_M1_CDNS_2 $T=98120 140130 0 0 $X=98040 $Y=139880
X155 1 M2_M1_CDNS_2 $T=98120 141740 0 0 $X=98040 $Y=141490
X156 1 M2_M1_CDNS_2 $T=98120 213330 0 0 $X=98040 $Y=213080
X157 1 M2_M1_CDNS_2 $T=98120 214940 0 0 $X=98040 $Y=214690
X158 1 M2_M1_CDNS_2 $T=98120 286530 0 0 $X=98040 $Y=286280
X159 1 M2_M1_CDNS_2 $T=98120 288140 0 0 $X=98040 $Y=287890
X160 2 M2_M1_CDNS_2 $T=112510 72600 0 0 $X=112430 $Y=72350
X161 2 M2_M1_CDNS_2 $T=112510 145800 0 0 $X=112430 $Y=145550
X162 2 M2_M1_CDNS_2 $T=112510 219000 0 0 $X=112430 $Y=218750
X163 15 M2_M1_CDNS_2 $T=112670 60970 0 0 $X=112590 $Y=60720
X164 16 M2_M1_CDNS_2 $T=112670 134170 0 0 $X=112590 $Y=133920
X165 17 M2_M1_CDNS_2 $T=112670 207370 0 0 $X=112590 $Y=207120
X166 18 M2_M1_CDNS_2 $T=112700 60050 0 0 $X=112620 $Y=59800
X167 19 M2_M1_CDNS_2 $T=112700 133250 0 0 $X=112620 $Y=133000
X168 20 M2_M1_CDNS_2 $T=112700 206450 0 0 $X=112620 $Y=206200
X169 21 M2_M1_CDNS_2 $T=112730 59100 0 0 $X=112650 $Y=58850
X170 22 M2_M1_CDNS_2 $T=112730 132300 0 0 $X=112650 $Y=132050
X171 23 M2_M1_CDNS_2 $T=112730 205500 0 0 $X=112650 $Y=205250
X172 24 M2_M1_CDNS_2 $T=112800 65320 0 0 $X=112720 $Y=65070
X173 25 M2_M1_CDNS_2 $T=112800 138520 0 0 $X=112720 $Y=138270
X174 26 M2_M1_CDNS_2 $T=112800 211720 0 0 $X=112720 $Y=211470
X175 27 M2_M1_CDNS_2 $T=114770 6460 0 0 $X=114690 $Y=6210
X176 28 M2_M1_CDNS_2 $T=114770 79660 0 0 $X=114690 $Y=79410
X177 29 M2_M1_CDNS_2 $T=114770 152860 0 0 $X=114690 $Y=152610
X178 30 M2_M1_CDNS_2 $T=114770 226060 0 0 $X=114690 $Y=225810
X179 1 M2_M1_CDNS_2 $T=125760 68120 0 0 $X=125680 $Y=67870
X180 1 M2_M1_CDNS_2 $T=125760 141320 0 0 $X=125680 $Y=141070
X181 1 M2_M1_CDNS_2 $T=125760 214520 0 0 $X=125680 $Y=214270
X182 1 M2_M1_CDNS_2 $T=127790 68120 0 0 $X=127710 $Y=67870
X183 1 M2_M1_CDNS_2 $T=127790 141320 0 0 $X=127710 $Y=141070
X184 1 M2_M1_CDNS_2 $T=127790 214520 0 0 $X=127710 $Y=214270
X185 15 M2_M1_CDNS_2 $T=127930 57970 0 0 $X=127850 $Y=57720
X186 16 M2_M1_CDNS_2 $T=127930 131170 0 0 $X=127850 $Y=130920
X187 17 M2_M1_CDNS_2 $T=127930 204370 0 0 $X=127850 $Y=204120
X188 18 M2_M1_CDNS_2 $T=128370 60020 0 0 $X=128290 $Y=59770
X189 19 M2_M1_CDNS_2 $T=128370 133220 0 0 $X=128290 $Y=132970
X190 20 M2_M1_CDNS_2 $T=128370 206420 0 0 $X=128290 $Y=206170
X191 1 M2_M1_CDNS_2 $T=162210 66930 0 0 $X=162130 $Y=66680
X192 1 M2_M1_CDNS_2 $T=162210 68540 0 0 $X=162130 $Y=68290
X193 1 M2_M1_CDNS_2 $T=162210 140130 0 0 $X=162130 $Y=139880
X194 1 M2_M1_CDNS_2 $T=162210 141740 0 0 $X=162130 $Y=141490
X195 1 M2_M1_CDNS_2 $T=162210 213330 0 0 $X=162130 $Y=213080
X196 1 M2_M1_CDNS_2 $T=162210 214940 0 0 $X=162130 $Y=214690
X197 1 M2_M1_CDNS_2 $T=162210 286530 0 0 $X=162130 $Y=286280
X198 1 M2_M1_CDNS_2 $T=162210 288140 0 0 $X=162130 $Y=287890
X199 2 M2_M1_CDNS_2 $T=176600 72600 0 0 $X=176520 $Y=72350
X200 2 M2_M1_CDNS_2 $T=176600 145800 0 0 $X=176520 $Y=145550
X201 2 M2_M1_CDNS_2 $T=176600 219000 0 0 $X=176520 $Y=218750
X202 31 M2_M1_CDNS_2 $T=176760 60970 0 0 $X=176680 $Y=60720
X203 32 M2_M1_CDNS_2 $T=176760 134170 0 0 $X=176680 $Y=133920
X204 33 M2_M1_CDNS_2 $T=176760 207370 0 0 $X=176680 $Y=207120
X205 34 M2_M1_CDNS_2 $T=176790 60050 0 0 $X=176710 $Y=59800
X206 35 M2_M1_CDNS_2 $T=176790 133250 0 0 $X=176710 $Y=133000
X207 36 M2_M1_CDNS_2 $T=176790 206450 0 0 $X=176710 $Y=206200
X208 37 M2_M1_CDNS_2 $T=176820 59100 0 0 $X=176740 $Y=58850
X209 38 M2_M1_CDNS_2 $T=176820 132300 0 0 $X=176740 $Y=132050
X210 39 M2_M1_CDNS_2 $T=176820 205500 0 0 $X=176740 $Y=205250
X211 40 M2_M1_CDNS_2 $T=176890 65320 0 0 $X=176810 $Y=65070
X212 41 M2_M1_CDNS_2 $T=176890 138520 0 0 $X=176810 $Y=138270
X213 42 M2_M1_CDNS_2 $T=176890 211720 0 0 $X=176810 $Y=211470
X214 43 M2_M1_CDNS_2 $T=178860 6460 0 0 $X=178780 $Y=6210
X215 44 M2_M1_CDNS_2 $T=178860 79660 0 0 $X=178780 $Y=79410
X216 45 M2_M1_CDNS_2 $T=178860 152860 0 0 $X=178780 $Y=152610
X217 46 M2_M1_CDNS_2 $T=178860 226060 0 0 $X=178780 $Y=225810
X218 1 M2_M1_CDNS_2 $T=189850 68120 0 0 $X=189770 $Y=67870
X219 1 M2_M1_CDNS_2 $T=189850 141320 0 0 $X=189770 $Y=141070
X220 1 M2_M1_CDNS_2 $T=189850 214520 0 0 $X=189770 $Y=214270
X221 1 M2_M1_CDNS_2 $T=191880 68120 0 0 $X=191800 $Y=67870
X222 1 M2_M1_CDNS_2 $T=191880 141320 0 0 $X=191800 $Y=141070
X223 1 M2_M1_CDNS_2 $T=191880 214520 0 0 $X=191800 $Y=214270
X224 31 M2_M1_CDNS_2 $T=192020 57970 0 0 $X=191940 $Y=57720
X225 32 M2_M1_CDNS_2 $T=192020 131170 0 0 $X=191940 $Y=130920
X226 33 M2_M1_CDNS_2 $T=192020 204370 0 0 $X=191940 $Y=204120
X227 34 M2_M1_CDNS_2 $T=192460 60020 0 0 $X=192380 $Y=59770
X228 35 M2_M1_CDNS_2 $T=192460 133220 0 0 $X=192380 $Y=132970
X229 36 M2_M1_CDNS_2 $T=192460 206420 0 0 $X=192380 $Y=206170
X230 47 M2_M1_CDNS_2 $T=242950 6460 0 0 $X=242870 $Y=6210
X231 48 M2_M1_CDNS_2 $T=242950 79660 0 0 $X=242870 $Y=79410
X232 49 M2_M1_CDNS_2 $T=242950 152860 0 0 $X=242870 $Y=152610
X233 50 M2_M1_CDNS_2 $T=242950 226060 0 0 $X=242870 $Y=225810
X234 3 M4_M3_CDNS_3 $T=41890 60920 0 0 $X=41810 $Y=60670
X235 4 M4_M3_CDNS_3 $T=41890 134120 0 0 $X=41810 $Y=133870
X236 5 M4_M3_CDNS_3 $T=41890 207320 0 0 $X=41810 $Y=207070
X237 51 M4_M3_CDNS_3 $T=41890 280520 0 0 $X=41810 $Y=280270
X238 9 M4_M3_CDNS_3 $T=42070 59420 0 0 $X=41990 $Y=59170
X239 10 M4_M3_CDNS_3 $T=42070 132620 0 0 $X=41990 $Y=132370
X240 11 M4_M3_CDNS_3 $T=42070 205820 0 0 $X=41990 $Y=205570
X241 9 M4_M3_CDNS_3 $T=75190 57370 0 90 $X=74940 $Y=57290
X242 10 M4_M3_CDNS_3 $T=75190 130570 0 90 $X=74940 $Y=130490
X243 11 M4_M3_CDNS_3 $T=75190 203770 0 90 $X=74940 $Y=203690
X244 52 M4_M3_CDNS_3 $T=75190 276970 0 90 $X=74940 $Y=276890
X245 6 M4_M3_CDNS_3 $T=93040 57940 0 0 $X=92960 $Y=57690
X246 7 M4_M3_CDNS_3 $T=93040 131140 0 0 $X=92960 $Y=130890
X247 8 M4_M3_CDNS_3 $T=93040 204340 0 0 $X=92960 $Y=204090
X248 53 M4_M3_CDNS_3 $T=93040 277540 0 0 $X=92960 $Y=277290
X249 15 M4_M3_CDNS_3 $T=105980 60920 0 0 $X=105900 $Y=60670
X250 16 M4_M3_CDNS_3 $T=105980 134120 0 0 $X=105900 $Y=133870
X251 17 M4_M3_CDNS_3 $T=105980 207320 0 0 $X=105900 $Y=207070
X252 54 M4_M3_CDNS_3 $T=105980 280520 0 0 $X=105900 $Y=280270
X253 21 M4_M3_CDNS_3 $T=106160 59420 0 0 $X=106080 $Y=59170
X254 22 M4_M3_CDNS_3 $T=106160 132620 0 0 $X=106080 $Y=132370
X255 23 M4_M3_CDNS_3 $T=106160 205820 0 0 $X=106080 $Y=205570
X256 21 M4_M3_CDNS_3 $T=139280 57370 0 90 $X=139030 $Y=57290
X257 22 M4_M3_CDNS_3 $T=139280 130570 0 90 $X=139030 $Y=130490
X258 23 M4_M3_CDNS_3 $T=139280 203770 0 90 $X=139030 $Y=203690
X259 55 M4_M3_CDNS_3 $T=139280 276970 0 90 $X=139030 $Y=276890
X260 18 M4_M3_CDNS_3 $T=157130 57940 0 0 $X=157050 $Y=57690
X261 19 M4_M3_CDNS_3 $T=157130 131140 0 0 $X=157050 $Y=130890
X262 20 M4_M3_CDNS_3 $T=157130 204340 0 0 $X=157050 $Y=204090
X263 56 M4_M3_CDNS_3 $T=157130 277540 0 0 $X=157050 $Y=277290
X264 31 M4_M3_CDNS_3 $T=170070 60920 0 0 $X=169990 $Y=60670
X265 32 M4_M3_CDNS_3 $T=170070 134120 0 0 $X=169990 $Y=133870
X266 33 M4_M3_CDNS_3 $T=170070 207320 0 0 $X=169990 $Y=207070
X267 57 M4_M3_CDNS_3 $T=170070 280520 0 0 $X=169990 $Y=280270
X268 37 M4_M3_CDNS_3 $T=170250 59420 0 0 $X=170170 $Y=59170
X269 38 M4_M3_CDNS_3 $T=170250 132620 0 0 $X=170170 $Y=132370
X270 39 M4_M3_CDNS_3 $T=170250 205820 0 0 $X=170170 $Y=205570
X271 37 M4_M3_CDNS_3 $T=203370 57370 0 90 $X=203120 $Y=57290
X272 38 M4_M3_CDNS_3 $T=203370 130570 0 90 $X=203120 $Y=130490
X273 39 M4_M3_CDNS_3 $T=203370 203770 0 90 $X=203120 $Y=203690
X274 58 M4_M3_CDNS_3 $T=203370 276970 0 90 $X=203120 $Y=276890
X275 34 M4_M3_CDNS_3 $T=221220 57940 0 0 $X=221140 $Y=57690
X276 35 M4_M3_CDNS_3 $T=221220 131140 0 0 $X=221140 $Y=130890
X277 36 M4_M3_CDNS_3 $T=221220 204340 0 0 $X=221140 $Y=204090
X278 59 M4_M3_CDNS_3 $T=221220 277540 0 0 $X=221140 $Y=277290
X279 2 M3_M2_CDNS_4 $T=38010 72260 0 0 $X=37930 $Y=72130
X280 2 M3_M2_CDNS_4 $T=38010 145460 0 0 $X=37930 $Y=145330
X281 2 M3_M2_CDNS_4 $T=38010 218660 0 0 $X=37930 $Y=218530
X282 6 M3_M2_CDNS_4 $T=46770 60050 0 0 $X=46690 $Y=59920
X283 7 M3_M2_CDNS_4 $T=46770 133250 0 0 $X=46690 $Y=133120
X284 8 M3_M2_CDNS_4 $T=46770 206450 0 0 $X=46690 $Y=206320
X285 27 M3_M2_CDNS_4 $T=57900 1030 0 0 $X=57820 $Y=900
X286 28 M3_M2_CDNS_4 $T=57900 74230 0 0 $X=57820 $Y=74100
X287 29 M3_M2_CDNS_4 $T=57900 147430 0 0 $X=57820 $Y=147300
X288 30 M3_M2_CDNS_4 $T=57900 220630 0 0 $X=57820 $Y=220500
X289 9 M3_M2_CDNS_4 $T=64230 55260 0 0 $X=64150 $Y=55130
X290 10 M3_M2_CDNS_4 $T=64230 128460 0 0 $X=64150 $Y=128330
X291 11 M3_M2_CDNS_4 $T=64230 201660 0 0 $X=64150 $Y=201530
X292 52 M3_M2_CDNS_4 $T=64230 274860 0 0 $X=64150 $Y=274730
X293 53 M3_M2_CDNS_4 $T=64280 279630 0 0 $X=64200 $Y=279500
X294 3 M3_M2_CDNS_4 $T=66720 57280 0 90 $X=66590 $Y=57200
X295 4 M3_M2_CDNS_4 $T=66720 130480 0 90 $X=66590 $Y=130400
X296 5 M3_M2_CDNS_4 $T=66720 203680 0 90 $X=66590 $Y=203600
X297 51 M3_M2_CDNS_4 $T=66720 276880 0 90 $X=66590 $Y=276800
X298 2 M3_M2_CDNS_4 $T=102100 72260 0 0 $X=102020 $Y=72130
X299 2 M3_M2_CDNS_4 $T=102100 145460 0 0 $X=102020 $Y=145330
X300 2 M3_M2_CDNS_4 $T=102100 218660 0 0 $X=102020 $Y=218530
X301 18 M3_M2_CDNS_4 $T=110860 60050 0 0 $X=110780 $Y=59920
X302 19 M3_M2_CDNS_4 $T=110860 133250 0 0 $X=110780 $Y=133120
X303 20 M3_M2_CDNS_4 $T=110860 206450 0 0 $X=110780 $Y=206320
X304 43 M3_M2_CDNS_4 $T=121990 1030 0 0 $X=121910 $Y=900
X305 44 M3_M2_CDNS_4 $T=121990 74230 0 0 $X=121910 $Y=74100
X306 45 M3_M2_CDNS_4 $T=121990 147430 0 0 $X=121910 $Y=147300
X307 46 M3_M2_CDNS_4 $T=121990 220630 0 0 $X=121910 $Y=220500
X308 21 M3_M2_CDNS_4 $T=128320 55260 0 0 $X=128240 $Y=55130
X309 22 M3_M2_CDNS_4 $T=128320 128460 0 0 $X=128240 $Y=128330
X310 23 M3_M2_CDNS_4 $T=128320 201660 0 0 $X=128240 $Y=201530
X311 55 M3_M2_CDNS_4 $T=128320 274860 0 0 $X=128240 $Y=274730
X312 56 M3_M2_CDNS_4 $T=128370 279630 0 0 $X=128290 $Y=279500
X313 15 M3_M2_CDNS_4 $T=130810 57280 0 90 $X=130680 $Y=57200
X314 16 M3_M2_CDNS_4 $T=130810 130480 0 90 $X=130680 $Y=130400
X315 17 M3_M2_CDNS_4 $T=130810 203680 0 90 $X=130680 $Y=203600
X316 54 M3_M2_CDNS_4 $T=130810 276880 0 90 $X=130680 $Y=276800
X317 2 M3_M2_CDNS_4 $T=166190 72260 0 0 $X=166110 $Y=72130
X318 2 M3_M2_CDNS_4 $T=166190 145460 0 0 $X=166110 $Y=145330
X319 2 M3_M2_CDNS_4 $T=166190 218660 0 0 $X=166110 $Y=218530
X320 34 M3_M2_CDNS_4 $T=174950 60050 0 0 $X=174870 $Y=59920
X321 35 M3_M2_CDNS_4 $T=174950 133250 0 0 $X=174870 $Y=133120
X322 36 M3_M2_CDNS_4 $T=174950 206450 0 0 $X=174870 $Y=206320
X323 47 M3_M2_CDNS_4 $T=186080 1030 0 0 $X=186000 $Y=900
X324 48 M3_M2_CDNS_4 $T=186080 74230 0 0 $X=186000 $Y=74100
X325 49 M3_M2_CDNS_4 $T=186080 147430 0 0 $X=186000 $Y=147300
X326 50 M3_M2_CDNS_4 $T=186080 220630 0 0 $X=186000 $Y=220500
X327 37 M3_M2_CDNS_4 $T=192410 55260 0 0 $X=192330 $Y=55130
X328 38 M3_M2_CDNS_4 $T=192410 128460 0 0 $X=192330 $Y=128330
X329 39 M3_M2_CDNS_4 $T=192410 201660 0 0 $X=192330 $Y=201530
X330 58 M3_M2_CDNS_4 $T=192410 274860 0 0 $X=192330 $Y=274730
X331 59 M3_M2_CDNS_4 $T=192460 279630 0 0 $X=192380 $Y=279500
X332 31 M3_M2_CDNS_4 $T=194900 57280 0 90 $X=194770 $Y=57200
X333 32 M3_M2_CDNS_4 $T=194900 130480 0 90 $X=194770 $Y=130400
X334 33 M3_M2_CDNS_4 $T=194900 203680 0 90 $X=194770 $Y=203600
X335 57 M3_M2_CDNS_4 $T=194900 276880 0 90 $X=194770 $Y=276800
X336 12 M5_M4_CDNS_5 $T=14800 59980 0 0 $X=14720 $Y=59730
X337 13 M5_M4_CDNS_5 $T=14800 133180 0 0 $X=14720 $Y=132930
X338 14 M5_M4_CDNS_5 $T=14800 206380 0 0 $X=14720 $Y=206130
X339 60 M5_M4_CDNS_5 $T=14800 279580 0 0 $X=14720 $Y=279330
X340 9 M5_M4_CDNS_5 $T=31930 59320 0 0 $X=31850 $Y=59070
X341 10 M5_M4_CDNS_5 $T=31930 132520 0 0 $X=31850 $Y=132270
X342 11 M5_M4_CDNS_5 $T=31930 205720 0 0 $X=31850 $Y=205470
X343 52 M5_M4_CDNS_5 $T=31930 278920 0 0 $X=31850 $Y=278670
X344 51 M5_M4_CDNS_5 $T=41890 280520 0 0 $X=41810 $Y=280270
X345 12 M5_M4_CDNS_5 $T=42050 65680 0 0 $X=41970 $Y=65430
X346 13 M5_M4_CDNS_5 $T=42050 138880 0 0 $X=41970 $Y=138630
X347 14 M5_M4_CDNS_5 $T=42050 212080 0 0 $X=41970 $Y=211830
X348 60 M5_M4_CDNS_5 $T=42050 285280 0 0 $X=41970 $Y=285030
X349 52 M5_M4_CDNS_5 $T=42070 279020 0 0 $X=41990 $Y=278770
X350 12 M5_M4_CDNS_5 $T=65300 57480 0 0 $X=65220 $Y=57230
X351 13 M5_M4_CDNS_5 $T=65300 130680 0 0 $X=65220 $Y=130430
X352 14 M5_M4_CDNS_5 $T=65300 203880 0 0 $X=65220 $Y=203630
X353 60 M5_M4_CDNS_5 $T=65300 277080 0 0 $X=65220 $Y=276830
X354 9 M5_M4_CDNS_5 $T=75190 57370 0 90 $X=74940 $Y=57290
X355 10 M5_M4_CDNS_5 $T=75190 130570 0 90 $X=74940 $Y=130490
X356 11 M5_M4_CDNS_5 $T=75190 203770 0 90 $X=74940 $Y=203690
X357 52 M5_M4_CDNS_5 $T=75190 276970 0 90 $X=74940 $Y=276890
X358 24 M5_M4_CDNS_5 $T=78890 59980 0 0 $X=78810 $Y=59730
X359 25 M5_M4_CDNS_5 $T=78890 133180 0 0 $X=78810 $Y=132930
X360 26 M5_M4_CDNS_5 $T=78890 206380 0 0 $X=78810 $Y=206130
X361 61 M5_M4_CDNS_5 $T=78890 279580 0 0 $X=78810 $Y=279330
X362 3 M5_M4_CDNS_5 $T=84220 57420 0 0 $X=84140 $Y=57170
X363 4 M5_M4_CDNS_5 $T=84220 130620 0 0 $X=84140 $Y=130370
X364 5 M5_M4_CDNS_5 $T=84220 203820 0 0 $X=84140 $Y=203570
X365 51 M5_M4_CDNS_5 $T=84220 277020 0 0 $X=84140 $Y=276770
X366 6 M5_M4_CDNS_5 $T=93040 57940 0 0 $X=92960 $Y=57690
X367 7 M5_M4_CDNS_5 $T=93040 131140 0 0 $X=92960 $Y=130890
X368 8 M5_M4_CDNS_5 $T=93040 204340 0 0 $X=92960 $Y=204090
X369 53 M5_M4_CDNS_5 $T=93040 277540 0 0 $X=92960 $Y=277290
X370 21 M5_M4_CDNS_5 $T=96020 59320 0 0 $X=95940 $Y=59070
X371 22 M5_M4_CDNS_5 $T=96020 132520 0 0 $X=95940 $Y=132270
X372 23 M5_M4_CDNS_5 $T=96020 205720 0 0 $X=95940 $Y=205470
X373 55 M5_M4_CDNS_5 $T=96020 278920 0 0 $X=95940 $Y=278670
X374 54 M5_M4_CDNS_5 $T=105980 280520 0 0 $X=105900 $Y=280270
X375 24 M5_M4_CDNS_5 $T=106140 65680 0 0 $X=106060 $Y=65430
X376 25 M5_M4_CDNS_5 $T=106140 138880 0 0 $X=106060 $Y=138630
X377 26 M5_M4_CDNS_5 $T=106140 212080 0 0 $X=106060 $Y=211830
X378 61 M5_M4_CDNS_5 $T=106140 285280 0 0 $X=106060 $Y=285030
X379 55 M5_M4_CDNS_5 $T=106160 279020 0 0 $X=106080 $Y=278770
X380 24 M5_M4_CDNS_5 $T=129390 57480 0 0 $X=129310 $Y=57230
X381 25 M5_M4_CDNS_5 $T=129390 130680 0 0 $X=129310 $Y=130430
X382 26 M5_M4_CDNS_5 $T=129390 203880 0 0 $X=129310 $Y=203630
X383 61 M5_M4_CDNS_5 $T=129390 277080 0 0 $X=129310 $Y=276830
X384 21 M5_M4_CDNS_5 $T=139280 57370 0 90 $X=139030 $Y=57290
X385 22 M5_M4_CDNS_5 $T=139280 130570 0 90 $X=139030 $Y=130490
X386 23 M5_M4_CDNS_5 $T=139280 203770 0 90 $X=139030 $Y=203690
X387 55 M5_M4_CDNS_5 $T=139280 276970 0 90 $X=139030 $Y=276890
X388 40 M5_M4_CDNS_5 $T=142980 59980 0 0 $X=142900 $Y=59730
X389 41 M5_M4_CDNS_5 $T=142980 133180 0 0 $X=142900 $Y=132930
X390 42 M5_M4_CDNS_5 $T=142980 206380 0 0 $X=142900 $Y=206130
X391 62 M5_M4_CDNS_5 $T=142980 279580 0 0 $X=142900 $Y=279330
X392 15 M5_M4_CDNS_5 $T=148310 57420 0 0 $X=148230 $Y=57170
X393 16 M5_M4_CDNS_5 $T=148310 130620 0 0 $X=148230 $Y=130370
X394 17 M5_M4_CDNS_5 $T=148310 203820 0 0 $X=148230 $Y=203570
X395 54 M5_M4_CDNS_5 $T=148310 277020 0 0 $X=148230 $Y=276770
X396 18 M5_M4_CDNS_5 $T=157130 57940 0 0 $X=157050 $Y=57690
X397 19 M5_M4_CDNS_5 $T=157130 131140 0 0 $X=157050 $Y=130890
X398 20 M5_M4_CDNS_5 $T=157130 204340 0 0 $X=157050 $Y=204090
X399 56 M5_M4_CDNS_5 $T=157130 277540 0 0 $X=157050 $Y=277290
X400 37 M5_M4_CDNS_5 $T=160110 59320 0 0 $X=160030 $Y=59070
X401 38 M5_M4_CDNS_5 $T=160110 132520 0 0 $X=160030 $Y=132270
X402 39 M5_M4_CDNS_5 $T=160110 205720 0 0 $X=160030 $Y=205470
X403 58 M5_M4_CDNS_5 $T=160110 278920 0 0 $X=160030 $Y=278670
X404 57 M5_M4_CDNS_5 $T=170070 280520 0 0 $X=169990 $Y=280270
X405 40 M5_M4_CDNS_5 $T=170230 65680 0 0 $X=170150 $Y=65430
X406 41 M5_M4_CDNS_5 $T=170230 138880 0 0 $X=170150 $Y=138630
X407 42 M5_M4_CDNS_5 $T=170230 212080 0 0 $X=170150 $Y=211830
X408 62 M5_M4_CDNS_5 $T=170230 285280 0 0 $X=170150 $Y=285030
X409 58 M5_M4_CDNS_5 $T=170250 279020 0 0 $X=170170 $Y=278770
X410 40 M5_M4_CDNS_5 $T=193480 57480 0 0 $X=193400 $Y=57230
X411 41 M5_M4_CDNS_5 $T=193480 130680 0 0 $X=193400 $Y=130430
X412 42 M5_M4_CDNS_5 $T=193480 203880 0 0 $X=193400 $Y=203630
X413 62 M5_M4_CDNS_5 $T=193480 277080 0 0 $X=193400 $Y=276830
X414 37 M5_M4_CDNS_5 $T=203370 57370 0 90 $X=203120 $Y=57290
X415 38 M5_M4_CDNS_5 $T=203370 130570 0 90 $X=203120 $Y=130490
X416 39 M5_M4_CDNS_5 $T=203370 203770 0 90 $X=203120 $Y=203690
X417 58 M5_M4_CDNS_5 $T=203370 276970 0 90 $X=203120 $Y=276890
X418 31 M5_M4_CDNS_5 $T=212400 57420 0 0 $X=212320 $Y=57170
X419 32 M5_M4_CDNS_5 $T=212400 130620 0 0 $X=212320 $Y=130370
X420 33 M5_M4_CDNS_5 $T=212400 203820 0 0 $X=212320 $Y=203570
X421 57 M5_M4_CDNS_5 $T=212400 277020 0 0 $X=212320 $Y=276770
X422 34 M5_M4_CDNS_5 $T=221220 57940 0 0 $X=221140 $Y=57690
X423 35 M5_M4_CDNS_5 $T=221220 131140 0 0 $X=221140 $Y=130890
X424 36 M5_M4_CDNS_5 $T=221220 204340 0 0 $X=221140 $Y=204090
X425 59 M5_M4_CDNS_5 $T=221220 277540 0 0 $X=221140 $Y=277290
X426 12 M4_M3_CDNS_6 $T=14800 59980 0 0 $X=14720 $Y=59730
X427 13 M4_M3_CDNS_6 $T=14800 133180 0 0 $X=14720 $Y=132930
X428 14 M4_M3_CDNS_6 $T=14800 206380 0 0 $X=14720 $Y=206130
X429 60 M4_M3_CDNS_6 $T=14800 279580 0 0 $X=14720 $Y=279330
X430 3 M4_M3_CDNS_6 $T=30970 60910 0 0 $X=30890 $Y=60660
X431 4 M4_M3_CDNS_6 $T=30970 134110 0 0 $X=30890 $Y=133860
X432 5 M4_M3_CDNS_6 $T=30970 207310 0 0 $X=30890 $Y=207060
X433 51 M4_M3_CDNS_6 $T=30970 280510 0 0 $X=30890 $Y=280260
X434 9 M4_M3_CDNS_6 $T=31930 59320 0 0 $X=31850 $Y=59070
X435 10 M4_M3_CDNS_6 $T=31930 132520 0 0 $X=31850 $Y=132270
X436 11 M4_M3_CDNS_6 $T=31930 205720 0 0 $X=31850 $Y=205470
X437 52 M4_M3_CDNS_6 $T=31930 278920 0 0 $X=31850 $Y=278670
X438 12 M4_M3_CDNS_6 $T=42050 65680 0 0 $X=41970 $Y=65430
X439 13 M4_M3_CDNS_6 $T=42050 138880 0 0 $X=41970 $Y=138630
X440 14 M4_M3_CDNS_6 $T=42050 212080 0 0 $X=41970 $Y=211830
X441 60 M4_M3_CDNS_6 $T=42050 285280 0 0 $X=41970 $Y=285030
X442 52 M4_M3_CDNS_6 $T=42070 279020 0 0 $X=41990 $Y=278770
X443 12 M4_M3_CDNS_6 $T=65300 57480 0 0 $X=65220 $Y=57230
X444 13 M4_M3_CDNS_6 $T=65300 130680 0 0 $X=65220 $Y=130430
X445 14 M4_M3_CDNS_6 $T=65300 203880 0 0 $X=65220 $Y=203630
X446 60 M4_M3_CDNS_6 $T=65300 277080 0 0 $X=65220 $Y=276830
X447 24 M4_M3_CDNS_6 $T=78890 59980 0 0 $X=78810 $Y=59730
X448 25 M4_M3_CDNS_6 $T=78890 133180 0 0 $X=78810 $Y=132930
X449 26 M4_M3_CDNS_6 $T=78890 206380 0 0 $X=78810 $Y=206130
X450 61 M4_M3_CDNS_6 $T=78890 279580 0 0 $X=78810 $Y=279330
X451 3 M4_M3_CDNS_6 $T=84220 57420 0 0 $X=84140 $Y=57170
X452 4 M4_M3_CDNS_6 $T=84220 130620 0 0 $X=84140 $Y=130370
X453 5 M4_M3_CDNS_6 $T=84220 203820 0 0 $X=84140 $Y=203570
X454 51 M4_M3_CDNS_6 $T=84220 277020 0 0 $X=84140 $Y=276770
X455 15 M4_M3_CDNS_6 $T=95060 60910 0 0 $X=94980 $Y=60660
X456 16 M4_M3_CDNS_6 $T=95060 134110 0 0 $X=94980 $Y=133860
X457 17 M4_M3_CDNS_6 $T=95060 207310 0 0 $X=94980 $Y=207060
X458 54 M4_M3_CDNS_6 $T=95060 280510 0 0 $X=94980 $Y=280260
X459 21 M4_M3_CDNS_6 $T=96020 59320 0 0 $X=95940 $Y=59070
X460 22 M4_M3_CDNS_6 $T=96020 132520 0 0 $X=95940 $Y=132270
X461 23 M4_M3_CDNS_6 $T=96020 205720 0 0 $X=95940 $Y=205470
X462 55 M4_M3_CDNS_6 $T=96020 278920 0 0 $X=95940 $Y=278670
X463 24 M4_M3_CDNS_6 $T=106140 65680 0 0 $X=106060 $Y=65430
X464 25 M4_M3_CDNS_6 $T=106140 138880 0 0 $X=106060 $Y=138630
X465 26 M4_M3_CDNS_6 $T=106140 212080 0 0 $X=106060 $Y=211830
X466 61 M4_M3_CDNS_6 $T=106140 285280 0 0 $X=106060 $Y=285030
X467 55 M4_M3_CDNS_6 $T=106160 279020 0 0 $X=106080 $Y=278770
X468 24 M4_M3_CDNS_6 $T=129390 57480 0 0 $X=129310 $Y=57230
X469 25 M4_M3_CDNS_6 $T=129390 130680 0 0 $X=129310 $Y=130430
X470 26 M4_M3_CDNS_6 $T=129390 203880 0 0 $X=129310 $Y=203630
X471 61 M4_M3_CDNS_6 $T=129390 277080 0 0 $X=129310 $Y=276830
X472 40 M4_M3_CDNS_6 $T=142980 59980 0 0 $X=142900 $Y=59730
X473 41 M4_M3_CDNS_6 $T=142980 133180 0 0 $X=142900 $Y=132930
X474 42 M4_M3_CDNS_6 $T=142980 206380 0 0 $X=142900 $Y=206130
X475 62 M4_M3_CDNS_6 $T=142980 279580 0 0 $X=142900 $Y=279330
X476 15 M4_M3_CDNS_6 $T=148310 57420 0 0 $X=148230 $Y=57170
X477 16 M4_M3_CDNS_6 $T=148310 130620 0 0 $X=148230 $Y=130370
X478 17 M4_M3_CDNS_6 $T=148310 203820 0 0 $X=148230 $Y=203570
X479 54 M4_M3_CDNS_6 $T=148310 277020 0 0 $X=148230 $Y=276770
X480 31 M4_M3_CDNS_6 $T=159150 60910 0 0 $X=159070 $Y=60660
X481 32 M4_M3_CDNS_6 $T=159150 134110 0 0 $X=159070 $Y=133860
X482 33 M4_M3_CDNS_6 $T=159150 207310 0 0 $X=159070 $Y=207060
X483 57 M4_M3_CDNS_6 $T=159150 280510 0 0 $X=159070 $Y=280260
X484 37 M4_M3_CDNS_6 $T=160110 59320 0 0 $X=160030 $Y=59070
X485 38 M4_M3_CDNS_6 $T=160110 132520 0 0 $X=160030 $Y=132270
X486 39 M4_M3_CDNS_6 $T=160110 205720 0 0 $X=160030 $Y=205470
X487 58 M4_M3_CDNS_6 $T=160110 278920 0 0 $X=160030 $Y=278670
X488 40 M4_M3_CDNS_6 $T=170230 65680 0 0 $X=170150 $Y=65430
X489 41 M4_M3_CDNS_6 $T=170230 138880 0 0 $X=170150 $Y=138630
X490 42 M4_M3_CDNS_6 $T=170230 212080 0 0 $X=170150 $Y=211830
X491 62 M4_M3_CDNS_6 $T=170230 285280 0 0 $X=170150 $Y=285030
X492 58 M4_M3_CDNS_6 $T=170250 279020 0 0 $X=170170 $Y=278770
X493 40 M4_M3_CDNS_6 $T=193480 57480 0 0 $X=193400 $Y=57230
X494 41 M4_M3_CDNS_6 $T=193480 130680 0 0 $X=193400 $Y=130430
X495 42 M4_M3_CDNS_6 $T=193480 203880 0 0 $X=193400 $Y=203630
X496 62 M4_M3_CDNS_6 $T=193480 277080 0 0 $X=193400 $Y=276830
X497 31 M4_M3_CDNS_6 $T=212400 57420 0 0 $X=212320 $Y=57170
X498 32 M4_M3_CDNS_6 $T=212400 130620 0 0 $X=212320 $Y=130370
X499 33 M4_M3_CDNS_6 $T=212400 203820 0 0 $X=212320 $Y=203570
X500 57 M4_M3_CDNS_6 $T=212400 277020 0 0 $X=212320 $Y=276770
X501 12 M3_M2_CDNS_7 $T=14800 59980 0 0 $X=14720 $Y=59730
X502 13 M3_M2_CDNS_7 $T=14800 133180 0 0 $X=14720 $Y=132930
X503 14 M3_M2_CDNS_7 $T=14800 206380 0 0 $X=14720 $Y=206130
X504 60 M3_M2_CDNS_7 $T=14800 279580 0 0 $X=14720 $Y=279330
X505 3 M3_M2_CDNS_7 $T=30970 60910 0 0 $X=30890 $Y=60660
X506 4 M3_M2_CDNS_7 $T=30970 134110 0 0 $X=30890 $Y=133860
X507 5 M3_M2_CDNS_7 $T=30970 207310 0 0 $X=30890 $Y=207060
X508 51 M3_M2_CDNS_7 $T=30970 280510 0 0 $X=30890 $Y=280260
X509 9 M3_M2_CDNS_7 $T=31930 59320 0 0 $X=31850 $Y=59070
X510 10 M3_M2_CDNS_7 $T=31930 132520 0 0 $X=31850 $Y=132270
X511 11 M3_M2_CDNS_7 $T=31930 205720 0 0 $X=31850 $Y=205470
X512 52 M3_M2_CDNS_7 $T=31930 278920 0 0 $X=31850 $Y=278670
X513 12 M3_M2_CDNS_7 $T=42050 65680 0 0 $X=41970 $Y=65430
X514 13 M3_M2_CDNS_7 $T=42050 138880 0 0 $X=41970 $Y=138630
X515 14 M3_M2_CDNS_7 $T=42050 212080 0 0 $X=41970 $Y=211830
X516 60 M3_M2_CDNS_7 $T=42050 285280 0 0 $X=41970 $Y=285030
X517 52 M3_M2_CDNS_7 $T=42070 279020 0 0 $X=41990 $Y=278770
X518 12 M3_M2_CDNS_7 $T=65300 57480 0 0 $X=65220 $Y=57230
X519 13 M3_M2_CDNS_7 $T=65300 130680 0 0 $X=65220 $Y=130430
X520 14 M3_M2_CDNS_7 $T=65300 203880 0 0 $X=65220 $Y=203630
X521 60 M3_M2_CDNS_7 $T=65300 277080 0 0 $X=65220 $Y=276830
X522 24 M3_M2_CDNS_7 $T=78890 59980 0 0 $X=78810 $Y=59730
X523 25 M3_M2_CDNS_7 $T=78890 133180 0 0 $X=78810 $Y=132930
X524 26 M3_M2_CDNS_7 $T=78890 206380 0 0 $X=78810 $Y=206130
X525 61 M3_M2_CDNS_7 $T=78890 279580 0 0 $X=78810 $Y=279330
X526 3 M3_M2_CDNS_7 $T=84220 57420 0 0 $X=84140 $Y=57170
X527 4 M3_M2_CDNS_7 $T=84220 130620 0 0 $X=84140 $Y=130370
X528 5 M3_M2_CDNS_7 $T=84220 203820 0 0 $X=84140 $Y=203570
X529 51 M3_M2_CDNS_7 $T=84220 277020 0 0 $X=84140 $Y=276770
X530 15 M3_M2_CDNS_7 $T=95060 60910 0 0 $X=94980 $Y=60660
X531 16 M3_M2_CDNS_7 $T=95060 134110 0 0 $X=94980 $Y=133860
X532 17 M3_M2_CDNS_7 $T=95060 207310 0 0 $X=94980 $Y=207060
X533 54 M3_M2_CDNS_7 $T=95060 280510 0 0 $X=94980 $Y=280260
X534 21 M3_M2_CDNS_7 $T=96020 59320 0 0 $X=95940 $Y=59070
X535 22 M3_M2_CDNS_7 $T=96020 132520 0 0 $X=95940 $Y=132270
X536 23 M3_M2_CDNS_7 $T=96020 205720 0 0 $X=95940 $Y=205470
X537 55 M3_M2_CDNS_7 $T=96020 278920 0 0 $X=95940 $Y=278670
X538 24 M3_M2_CDNS_7 $T=106140 65680 0 0 $X=106060 $Y=65430
X539 25 M3_M2_CDNS_7 $T=106140 138880 0 0 $X=106060 $Y=138630
X540 26 M3_M2_CDNS_7 $T=106140 212080 0 0 $X=106060 $Y=211830
X541 61 M3_M2_CDNS_7 $T=106140 285280 0 0 $X=106060 $Y=285030
X542 55 M3_M2_CDNS_7 $T=106160 279020 0 0 $X=106080 $Y=278770
X543 24 M3_M2_CDNS_7 $T=129390 57480 0 0 $X=129310 $Y=57230
X544 25 M3_M2_CDNS_7 $T=129390 130680 0 0 $X=129310 $Y=130430
X545 26 M3_M2_CDNS_7 $T=129390 203880 0 0 $X=129310 $Y=203630
X546 61 M3_M2_CDNS_7 $T=129390 277080 0 0 $X=129310 $Y=276830
X547 40 M3_M2_CDNS_7 $T=142980 59980 0 0 $X=142900 $Y=59730
X548 41 M3_M2_CDNS_7 $T=142980 133180 0 0 $X=142900 $Y=132930
X549 42 M3_M2_CDNS_7 $T=142980 206380 0 0 $X=142900 $Y=206130
X550 62 M3_M2_CDNS_7 $T=142980 279580 0 0 $X=142900 $Y=279330
X551 15 M3_M2_CDNS_7 $T=148310 57420 0 0 $X=148230 $Y=57170
X552 16 M3_M2_CDNS_7 $T=148310 130620 0 0 $X=148230 $Y=130370
X553 17 M3_M2_CDNS_7 $T=148310 203820 0 0 $X=148230 $Y=203570
X554 54 M3_M2_CDNS_7 $T=148310 277020 0 0 $X=148230 $Y=276770
X555 31 M3_M2_CDNS_7 $T=159150 60910 0 0 $X=159070 $Y=60660
X556 32 M3_M2_CDNS_7 $T=159150 134110 0 0 $X=159070 $Y=133860
X557 33 M3_M2_CDNS_7 $T=159150 207310 0 0 $X=159070 $Y=207060
X558 57 M3_M2_CDNS_7 $T=159150 280510 0 0 $X=159070 $Y=280260
X559 37 M3_M2_CDNS_7 $T=160110 59320 0 0 $X=160030 $Y=59070
X560 38 M3_M2_CDNS_7 $T=160110 132520 0 0 $X=160030 $Y=132270
X561 39 M3_M2_CDNS_7 $T=160110 205720 0 0 $X=160030 $Y=205470
X562 58 M3_M2_CDNS_7 $T=160110 278920 0 0 $X=160030 $Y=278670
X563 40 M3_M2_CDNS_7 $T=170230 65680 0 0 $X=170150 $Y=65430
X564 41 M3_M2_CDNS_7 $T=170230 138880 0 0 $X=170150 $Y=138630
X565 42 M3_M2_CDNS_7 $T=170230 212080 0 0 $X=170150 $Y=211830
X566 62 M3_M2_CDNS_7 $T=170230 285280 0 0 $X=170150 $Y=285030
X567 58 M3_M2_CDNS_7 $T=170250 279020 0 0 $X=170170 $Y=278770
X568 40 M3_M2_CDNS_7 $T=193480 57480 0 0 $X=193400 $Y=57230
X569 41 M3_M2_CDNS_7 $T=193480 130680 0 0 $X=193400 $Y=130430
X570 42 M3_M2_CDNS_7 $T=193480 203880 0 0 $X=193400 $Y=203630
X571 62 M3_M2_CDNS_7 $T=193480 277080 0 0 $X=193400 $Y=276830
X572 31 M3_M2_CDNS_7 $T=212400 57420 0 0 $X=212320 $Y=57170
X573 32 M3_M2_CDNS_7 $T=212400 130620 0 0 $X=212320 $Y=130370
X574 33 M3_M2_CDNS_7 $T=212400 203820 0 0 $X=212320 $Y=203570
X575 57 M3_M2_CDNS_7 $T=212400 277020 0 0 $X=212320 $Y=276770
X576 2 M2_M1_CDNS_8 $T=56170 72600 0 0 $X=56090 $Y=72470
X577 2 M2_M1_CDNS_8 $T=56170 145800 0 0 $X=56090 $Y=145670
X578 2 M2_M1_CDNS_8 $T=56170 219000 0 0 $X=56090 $Y=218870
X579 9 M2_M1_CDNS_8 $T=64180 56760 0 90 $X=64050 $Y=56680
X580 10 M2_M1_CDNS_8 $T=64180 129960 0 90 $X=64050 $Y=129880
X581 11 M2_M1_CDNS_8 $T=64180 203160 0 90 $X=64050 $Y=203080
X582 12 M2_M1_CDNS_8 $T=64650 65320 0 0 $X=64570 $Y=65190
X583 13 M2_M1_CDNS_8 $T=64650 138520 0 0 $X=64570 $Y=138390
X584 14 M2_M1_CDNS_8 $T=64650 211720 0 0 $X=64570 $Y=211590
X585 2 M2_M1_CDNS_8 $T=120260 72600 0 0 $X=120180 $Y=72470
X586 2 M2_M1_CDNS_8 $T=120260 145800 0 0 $X=120180 $Y=145670
X587 2 M2_M1_CDNS_8 $T=120260 219000 0 0 $X=120180 $Y=218870
X588 21 M2_M1_CDNS_8 $T=128270 56760 0 90 $X=128140 $Y=56680
X589 22 M2_M1_CDNS_8 $T=128270 129960 0 90 $X=128140 $Y=129880
X590 23 M2_M1_CDNS_8 $T=128270 203160 0 90 $X=128140 $Y=203080
X591 24 M2_M1_CDNS_8 $T=128740 65320 0 0 $X=128660 $Y=65190
X592 25 M2_M1_CDNS_8 $T=128740 138520 0 0 $X=128660 $Y=138390
X593 26 M2_M1_CDNS_8 $T=128740 211720 0 0 $X=128660 $Y=211590
X594 2 M2_M1_CDNS_8 $T=184350 72600 0 0 $X=184270 $Y=72470
X595 2 M2_M1_CDNS_8 $T=184350 145800 0 0 $X=184270 $Y=145670
X596 2 M2_M1_CDNS_8 $T=184350 219000 0 0 $X=184270 $Y=218870
X597 37 M2_M1_CDNS_8 $T=192360 56760 0 90 $X=192230 $Y=56680
X598 38 M2_M1_CDNS_8 $T=192360 129960 0 90 $X=192230 $Y=129880
X599 39 M2_M1_CDNS_8 $T=192360 203160 0 90 $X=192230 $Y=203080
X600 40 M2_M1_CDNS_8 $T=192830 65320 0 0 $X=192750 $Y=65190
X601 41 M2_M1_CDNS_8 $T=192830 138520 0 0 $X=192750 $Y=138390
X602 42 M2_M1_CDNS_8 $T=192830 211720 0 0 $X=192750 $Y=211590
X603 3 M2_M1_CDNS_9 $T=30970 60910 0 0 $X=30890 $Y=60660
X604 4 M2_M1_CDNS_9 $T=30970 134110 0 0 $X=30890 $Y=133860
X605 5 M2_M1_CDNS_9 $T=30970 207310 0 0 $X=30890 $Y=207060
X606 51 M2_M1_CDNS_9 $T=30970 280510 0 0 $X=30890 $Y=280260
X607 15 M2_M1_CDNS_9 $T=95060 60910 0 0 $X=94980 $Y=60660
X608 16 M2_M1_CDNS_9 $T=95060 134110 0 0 $X=94980 $Y=133860
X609 17 M2_M1_CDNS_9 $T=95060 207310 0 0 $X=94980 $Y=207060
X610 54 M2_M1_CDNS_9 $T=95060 280510 0 0 $X=94980 $Y=280260
X611 31 M2_M1_CDNS_9 $T=159150 60910 0 0 $X=159070 $Y=60660
X612 32 M2_M1_CDNS_9 $T=159150 134110 0 0 $X=159070 $Y=133860
X613 33 M2_M1_CDNS_9 $T=159150 207310 0 0 $X=159070 $Y=207060
X614 57 M2_M1_CDNS_9 $T=159150 280510 0 0 $X=159070 $Y=280260
X615 3 M5_M4_CDNS_10 $T=30970 60910 0 0 $X=30890 $Y=60780
X616 4 M5_M4_CDNS_10 $T=30970 134110 0 0 $X=30890 $Y=133980
X617 5 M5_M4_CDNS_10 $T=30970 207310 0 0 $X=30890 $Y=207180
X618 51 M5_M4_CDNS_10 $T=30970 280510 0 0 $X=30890 $Y=280380
X619 3 M5_M4_CDNS_10 $T=41890 60920 0 0 $X=41810 $Y=60790
X620 4 M5_M4_CDNS_10 $T=41890 134120 0 0 $X=41810 $Y=133990
X621 5 M5_M4_CDNS_10 $T=41890 207320 0 0 $X=41810 $Y=207190
X622 9 M5_M4_CDNS_10 $T=42070 59420 0 0 $X=41990 $Y=59290
X623 10 M5_M4_CDNS_10 $T=42070 132620 0 0 $X=41990 $Y=132490
X624 11 M5_M4_CDNS_10 $T=42070 205820 0 0 $X=41990 $Y=205690
X625 15 M5_M4_CDNS_10 $T=95060 60910 0 0 $X=94980 $Y=60780
X626 16 M5_M4_CDNS_10 $T=95060 134110 0 0 $X=94980 $Y=133980
X627 17 M5_M4_CDNS_10 $T=95060 207310 0 0 $X=94980 $Y=207180
X628 54 M5_M4_CDNS_10 $T=95060 280510 0 0 $X=94980 $Y=280380
X629 15 M5_M4_CDNS_10 $T=105980 60920 0 0 $X=105900 $Y=60790
X630 16 M5_M4_CDNS_10 $T=105980 134120 0 0 $X=105900 $Y=133990
X631 17 M5_M4_CDNS_10 $T=105980 207320 0 0 $X=105900 $Y=207190
X632 21 M5_M4_CDNS_10 $T=106160 59420 0 0 $X=106080 $Y=59290
X633 22 M5_M4_CDNS_10 $T=106160 132620 0 0 $X=106080 $Y=132490
X634 23 M5_M4_CDNS_10 $T=106160 205820 0 0 $X=106080 $Y=205690
X635 31 M5_M4_CDNS_10 $T=159150 60910 0 0 $X=159070 $Y=60780
X636 32 M5_M4_CDNS_10 $T=159150 134110 0 0 $X=159070 $Y=133980
X637 33 M5_M4_CDNS_10 $T=159150 207310 0 0 $X=159070 $Y=207180
X638 57 M5_M4_CDNS_10 $T=159150 280510 0 0 $X=159070 $Y=280380
X639 31 M5_M4_CDNS_10 $T=170070 60920 0 0 $X=169990 $Y=60790
X640 32 M5_M4_CDNS_10 $T=170070 134120 0 0 $X=169990 $Y=133990
X641 33 M5_M4_CDNS_10 $T=170070 207320 0 0 $X=169990 $Y=207190
X642 37 M5_M4_CDNS_10 $T=170250 59420 0 0 $X=170170 $Y=59290
X643 38 M5_M4_CDNS_10 $T=170250 132620 0 0 $X=170170 $Y=132490
X644 39 M5_M4_CDNS_10 $T=170250 205820 0 0 $X=170170 $Y=205690
X645 63 64 65 66 67 68 69 12 70 2
+ 1 71 72 73 13 74 75 76 14 77
+ 78 79 80 60 81 82 83 84 85 86
+ 87 88 89 90 9 91 10 92 11 93
+ 52 94 95 51 5 4 3 96 97 98
+ 99 100 6 7 8 53 101 102 103 104
+ 30 29 28 27 105 106 107 108 109 110
+ 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 1720 1710 1700 1722 1712 1702
+ 1721 1711 1701 1726 1716 1706 1725 1715 1705 1724
+ 1723 1714 1713 1704 1703 1717 1707 1697 1719 1709
+ 1699 1718 1708 1698 333 332 331 472 471 470
+ 319 318 317 330 329 328 ph2p3_Matrix_vector_Multiplication $T=-650 60 0 0 $X=-390 $Y=0
X646 12 13 14 60 125 3 69 24 126 2
+ 1 127 72 4 25 128 129 5 26 130
+ 131 51 132 61 133 134 135 136 137 9
+ 10 11 52 138 21 6 22 7 23 8
+ 55 53 139 54 17 16 15 140 141 142
+ 143 144 18 19 20 56 27 28 29 30
+ 46 45 44 43 145 146 147 148 149 150
+ 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 3222 3212 3202 3224 3214 3204
+ 3223 3213 3203 3228 3218 3208 3227 3217 3207 3226
+ 3225 3216 3215 3206 3205 3219 3209 3199 3221 3211
+ 3201 3220 3210 3200 1835 1834 1833 1974 1973 1972
+ 1821 1820 1819 1832 1831 1830 ph2p3_Matrix_vector_Multiplication $T=63440 60 0 0 $X=63700 $Y=0
X647 24 25 26 61 165 15 69 40 166 2
+ 1 167 72 16 41 168 169 17 42 170
+ 171 54 172 62 173 174 175 176 177 21
+ 22 23 55 178 37 18 38 19 39 20
+ 58 56 179 57 33 32 31 180 181 182
+ 183 184 34 35 36 59 43 44 45 46
+ 50 49 48 47 185 186 187 188 189 190
+ 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 4724 4714 4704 4726 4716 4706
+ 4725 4715 4705 4730 4720 4710 4729 4719 4709 4728
+ 4727 4718 4717 4708 4707 4721 4711 4701 4723 4713
+ 4703 4722 4712 4702 3337 3336 3335 3476 3475 3474
+ 3323 3322 3321 3334 3333 3332 ph2p3_Matrix_vector_Multiplication $T=127530 60 0 0 $X=127790 $Y=0
X648 40 41 42 62 205 31 69 206 207 2
+ 1 208 72 32 209 210 211 33 212 213
+ 214 57 215 216 217 218 219 220 221 37
+ 38 39 58 222 223 34 224 35 225 36
+ 226 59 227 228 229 230 231 232 233 234
+ 235 236 237 238 239 240 47 48 49 50
+ 241 242 243 244 245 246 247 248 249 250
+ 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 6226 6216 6206 6228 6218 6208
+ 6227 6217 6207 6232 6222 6212 6231 6221 6211 6230
+ 6229 6220 6219 6210 6209 6223 6213 6203 6225 6215
+ 6205 6224 6214 6204 4839 4838 4837 4978 4977 4976
+ 4825 4824 4823 4836 4835 4834 ph2p3_Matrix_vector_Multiplication $T=191620 60 0 0 $X=191880 $Y=0
.ends ph3_sytolic_array
